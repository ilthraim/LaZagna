
module top (input clk, input reset,input [351:0] top_inp, output [143:0] top_outp); 
 


 wire [207:0] inp_dbram1;
wire [159:0] outp_dbram1;

dbram_2048_40bit_module_2 dbram1 (.clk(clk),.reset(reset),.inp(inp_dbram1),.outp(outp_dbram1)); 


 wire [835:0] inp_sysarr1;
wire [447:0] outp_sysarr1;

systolic_array_4_fp16bit_2 sysarr1 (.clk(clk),.reset(reset),.inp(inp_sysarr1),.outp(outp_sysarr1)); 
wire [159:0] inp_interface_1; 
wire [835:0] outp_interface_1; 

interface_1 inst_interface_1(.clk(clk),.reset(reset),.inp(inp_interface_1),.outp(outp_interface_1)); 


 wire [1727:0] inp_dbram2;
wire [1439:0] outp_dbram2;

dbram_2048_60bit_module_12 dbram2 (.clk(clk),.reset(reset),.inp(inp_dbram2),.outp(outp_dbram2)); 
wire [895:0] inp_interface_2; 
wire [1727:0] outp_interface_2; 

interface_2 inst_interface_2(.clk(clk),.reset(reset),.inp(inp_interface_2),.outp(outp_interface_2)); 


 wire [1059:0] inp_dbram3;
wire [799:0] outp_dbram3;

dbram_4096_40bit_module_10 dbram3 (.clk(clk),.reset(reset),.inp(inp_dbram3),.outp(outp_dbram3)); 
wire [895:0] inp_interface_3; 
wire [1059:0] outp_interface_3; 

interface_3 inst_interface_3(.clk(clk),.reset(reset),.inp(inp_interface_3),.outp(outp_interface_3)); 


 wire [835:0] inp_sysarr2;
wire [447:0] outp_sysarr2;

systolic_array_4_fp16bit_2 sysarr2 (.clk(clk),.reset(reset),.inp(inp_sysarr2),.outp(outp_sysarr2)); 
wire [799:0] inp_interface_4; 
wire [835:0] outp_interface_4; 

interface_4 inst_interface_4(.clk(clk),.reset(reset),.inp(inp_interface_4),.outp(outp_interface_4)); 


 wire [835:0] inp_sysarr3;
wire [447:0] outp_sysarr3;

systolic_array_4_fp16bit_2 sysarr3 (.clk(clk),.reset(reset),.inp(inp_sysarr3),.outp(outp_sysarr3)); 
wire [1439:0] inp_interface_5; 
wire [835:0] outp_interface_5; 

interface_5 inst_interface_5(.clk(clk),.reset(reset),.inp(inp_interface_5),.outp(outp_interface_5)); 


 wire [2919:0] inp_dbram4;
wire [2399:0] outp_dbram4;

dbram_4096_60bit_module_20 dbram4 (.clk(clk),.reset(reset),.inp(inp_dbram4),.outp(outp_dbram4)); 
wire [895:0] inp_interface_6; 
wire [2919:0] outp_interface_6; 

interface_6 inst_interface_6(.clk(clk),.reset(reset),.inp(inp_interface_6),.outp(outp_interface_6)); 


 wire [3095:0] inp_activ1;
wire [3083:0] outp_activ1;

activation_32_16bit_module_6 activ1 (.clk(clk),.reset(reset),.inp(inp_activ1),.outp(outp_activ1)); 
wire [2399:0] inp_interface_7; 
wire [3095:0] outp_interface_7; 

interface_7 inst_interface_7(.clk(clk),.reset(reset),.inp(inp_interface_7),.outp(outp_interface_7)); 


 wire [3131:0] inp_activ2;
wire [3095:0] outp_activ2;

activation_32_8bit_module_12 activ2 (.clk(clk),.reset(reset),.inp(inp_activ2),.outp(outp_activ2)); 
wire [2399:0] inp_interface_8; 
wire [3131:0] outp_interface_8; 

interface_8 inst_interface_8(.clk(clk),.reset(reset),.inp(inp_interface_8),.outp(outp_interface_8)); 


 wire [895:0] inp_adder_tree1;
wire [223:0] outp_adder_tree1;

adder_tree_3_8bit_14 adder_tree1 (.clk(clk),.reset(reset),.inp(inp_adder_tree1),.outp(outp_adder_tree1)); 
wire [1247:0] inp_interface_9; 
wire [895:0] outp_interface_9; 

interface_9 inst_interface_9(.clk(clk),.reset(reset),.inp(inp_interface_9),.outp(outp_interface_9)); 


 wire [1535:0] inp_adder_tree2;
wire [191:0] outp_adder_tree2;

adder_tree_4_4bit_24 adder_tree2 (.clk(clk),.reset(reset),.inp(inp_adder_tree2),.outp(outp_adder_tree2)); 
wire [1887:0] inp_interface_10; 
wire [1535:0] outp_interface_10; 

interface_10 inst_interface_10(.clk(clk),.reset(reset),.inp(inp_interface_10),.outp(outp_interface_10)); 


 wire [5119:0] inp_adder_tree3;
wire [639:0] outp_adder_tree3;

adder_tree_4_16bit_20 adder_tree3 (.clk(clk),.reset(reset),.inp(inp_adder_tree3),.outp(outp_adder_tree3)); 
wire [6595:0] inp_interface_11; 
wire [5119:0] outp_interface_11; 

interface_11 inst_interface_11(.clk(clk),.reset(reset),.inp(inp_interface_11),.outp(outp_interface_11)); 


 wire [835:0] inp_sysarr5;
wire [447:0] outp_sysarr5;

systolic_array_4_fp16bit_2 sysarr5 (.clk(clk),.reset(reset),.inp(inp_sysarr5),.outp(outp_sysarr5)); 
wire [6595:0] inp_interface_12; 
wire [835:0] outp_interface_12; 

interface_12 inst_interface_12(.clk(clk),.reset(reset),.inp(inp_interface_12),.outp(outp_interface_12)); 


 wire [143:0] inp_dbram5;
wire [119:0] outp_dbram5;

dbram_2048_60bit_module_1 dbram5 (.clk(clk),.reset(reset),.inp(inp_dbram5),.outp(outp_dbram5)); 


 wire [417:0] inp_sysarr4;
wire [223:0] outp_sysarr4;

systolic_array_4_fp16bit_1 sysarr4 (.clk(clk),.reset(reset),.inp(inp_sysarr4),.outp(outp_sysarr4)); 
wire [119:0] inp_interface_14; 
wire [417:0] outp_interface_14; 

interface_14 inst_interface_14(.clk(clk),.reset(reset),.inp(inp_interface_14),.outp(outp_interface_14)); 


 wire [127:0] inp_activ3;
wire [127:0] outp_activ3;

sigmoid_16bit_8 activ3 (.clk(clk),.reset(reset),.inp(inp_activ3),.outp(outp_activ3)); 
wire [223:0] inp_interface_15; 
wire [127:0] outp_interface_15; 

interface_15 inst_interface_15(.clk(clk),.reset(reset),.inp(inp_interface_15),.outp(outp_interface_15)); 


 wire [383:0] inp_adder_tree4;
wire [95:0] outp_adder_tree4;

adder_tree_3_8bit_6 adder_tree4 (.clk(clk),.reset(reset),.inp(inp_adder_tree4),.outp(outp_adder_tree4)); 
wire [119:0] inp_interface_16; 
wire [383:0] outp_interface_16; 

interface_16 inst_interface_16(.clk(clk),.reset(reset),.inp(inp_interface_16),.outp(outp_interface_16)); 


 wire [1151:0] inp_adder_tree5;
wire [143:0] outp_adder_tree5;

adder_tree_4_4bit_18 adder_tree5 (.clk(clk),.reset(reset),.inp(inp_adder_tree5),.outp(outp_adder_tree5)); 
wire [863:0] inp_interface_17; 
wire [1151:0] outp_interface_17; 

interface_17 inst_interface_17(.clk(clk),.reset(reset),.inp(inp_interface_17),.outp(outp_interface_17)); 

assign inp_dbram1 = top_inp[207:0]; 

assign inp_sysarr1 = outp_interface_1; 
assign inp_interface_1 = {outp_dbram1}; 
 

assign inp_dbram2 = outp_interface_2; 
assign inp_interface_2 = {outp_sysarr1,outp_sysarr5}; 
 

assign inp_dbram3 = outp_interface_3; 
assign inp_interface_3 = {outp_sysarr1,outp_sysarr5}; 
 

assign inp_sysarr2 = outp_interface_4; 
assign inp_interface_4 = {outp_dbram3}; 
 

assign inp_sysarr3 = outp_interface_5; 
assign inp_interface_5 = {outp_dbram2}; 
 

assign inp_dbram4 = outp_interface_6; 
assign inp_interface_6 = {outp_sysarr2,outp_sysarr3}; 
 

assign inp_activ1 = outp_interface_7; 
assign inp_interface_7 = {outp_dbram4}; 
 

assign inp_activ2 = outp_interface_8; 
assign inp_interface_8 = {outp_dbram4}; 
 

assign inp_adder_tree1 = outp_interface_9; 
assign inp_interface_9 = {outp_sysarr2,outp_dbram3}; 
 

assign inp_adder_tree2 = outp_interface_10; 
assign inp_interface_10 = {outp_sysarr3,outp_dbram2}; 
 

assign inp_adder_tree3 = outp_interface_11; 
assign inp_interface_11 = {outp_adder_tree1,outp_adder_tree2,outp_activ1,outp_activ2}; 
 

assign inp_sysarr5 = outp_interface_12; 
assign inp_interface_12 = {outp_adder_tree1,outp_adder_tree2,outp_activ1,outp_activ2}; 
 

assign inp_dbram5 = top_inp[351:208]; 

assign inp_sysarr4 = outp_interface_14; 
assign inp_interface_14 = {outp_dbram5}; 
 

assign inp_activ3 = outp_interface_15; 
assign inp_interface_15 = {outp_sysarr4}; 
 

assign inp_adder_tree4 = outp_interface_16; 
assign inp_interface_16 = {outp_dbram5}; 
 

assign inp_adder_tree5 = outp_interface_17; 
assign top_outp[143:0] = outp_adder_tree5; 
assign inp_interface_17 = {outp_activ3,outp_adder_tree4,outp_adder_tree3}; 
 

 endmodule 


module interface_1(input [159:0] inp, output reg [835:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[159:0] <= inp ; 
outp[319:160] <= inp ; 
outp[479:320] <= inp ; 
outp[639:480] <= inp ; 
outp[799:640] <= inp ; 
outp[835:800] <= inp[35:0] ; 
end 
endmodule 

module interface_2(input [895:0] inp, output reg [1727:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[895:0] <= inp ; 
outp[1727:896] <= inp[831:0] ; 
end 
endmodule 

module interface_3(input [895:0] inp, output reg [1059:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[895:0] <= inp ; 
outp[1059:896] <= inp[163:0] ; 
end 
endmodule 

module interface_4(input [799:0] inp, output reg [835:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[799:0] <= inp ; 
outp[835:800] <= inp[35:0] ; 
end 
endmodule 

module interface_5(input [1439:0] inp, output reg [835:0] outp, input clk, input reset);
reg [1439:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
wire [719:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
mux_module mux_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
xor_module xor_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
xor_module xor_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
mux_module mux_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
mux_module mux_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
mux_module mux_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
xor_module xor_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
mux_module mux_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
mux_module mux_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
xor_module xor_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
mux_module mux_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
xor_module xor_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
mux_module mux_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
xor_module xor_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
xor_module xor_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
xor_module xor_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
mux_module mux_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
xor_module xor_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
mux_module mux_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
mux_module mux_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
xor_module xor_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
mux_module mux_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
xor_module xor_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
mux_module mux_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
xor_module xor_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
mux_module mux_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
xor_module xor_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
xor_module xor_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
xor_module xor_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
mux_module mux_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
mux_module mux_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
xor_module xor_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
xor_module xor_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
mux_module mux_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
mux_module mux_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
xor_module xor_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
xor_module xor_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
xor_module xor_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
xor_module xor_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
xor_module xor_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
xor_module xor_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
mux_module mux_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
mux_module mux_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
xor_module xor_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
xor_module xor_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
xor_module xor_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
mux_module mux_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
mux_module mux_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
xor_module xor_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
mux_module mux_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
mux_module mux_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
xor_module xor_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
mux_module mux_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
mux_module mux_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
mux_module mux_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
mux_module mux_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
xor_module xor_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
mux_module mux_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
mux_module mux_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
xor_module xor_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
mux_module mux_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
xor_module xor_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
mux_module mux_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
mux_module mux_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
xor_module xor_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
xor_module xor_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
xor_module xor_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
xor_module xor_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
mux_module mux_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
xor_module xor_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
mux_module mux_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
mux_module mux_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
mux_module mux_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
mux_module mux_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
mux_module mux_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
xor_module xor_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
xor_module xor_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
xor_module xor_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
xor_module xor_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
mux_module mux_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
xor_module xor_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
mux_module mux_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
mux_module mux_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
mux_module mux_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
xor_module xor_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
xor_module xor_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
mux_module mux_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
xor_module xor_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
mux_module mux_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
xor_module xor_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
xor_module xor_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
xor_module xor_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
xor_module xor_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
xor_module xor_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
mux_module mux_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
mux_module mux_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
xor_module xor_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
xor_module xor_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
xor_module xor_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
xor_module xor_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
mux_module mux_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
xor_module xor_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
xor_module xor_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
mux_module mux_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
mux_module mux_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
xor_module xor_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
xor_module xor_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
xor_module xor_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
mux_module mux_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
xor_module xor_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
xor_module xor_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
xor_module xor_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
mux_module mux_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
xor_module xor_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
xor_module xor_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
mux_module mux_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
xor_module xor_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
mux_module mux_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
xor_module xor_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
xor_module xor_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
xor_module xor_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
mux_module mux_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
xor_module xor_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
mux_module mux_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
mux_module mux_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
xor_module xor_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
xor_module xor_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
mux_module mux_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
mux_module mux_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
mux_module mux_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
xor_module xor_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
xor_module xor_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
mux_module mux_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
mux_module mux_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
xor_module xor_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
xor_module xor_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
xor_module xor_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
xor_module xor_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
mux_module mux_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
mux_module mux_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
mux_module mux_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
xor_module xor_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
mux_module mux_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
xor_module xor_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
xor_module xor_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
mux_module mux_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
xor_module xor_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
mux_module mux_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
xor_module xor_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
xor_module xor_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
xor_module xor_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
mux_module mux_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
mux_module mux_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
xor_module xor_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
xor_module xor_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
mux_module mux_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
xor_module xor_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
mux_module mux_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
xor_module xor_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
mux_module mux_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
xor_module xor_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
mux_module mux_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
xor_module xor_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
xor_module xor_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
xor_module xor_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
mux_module mux_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
xor_module xor_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
mux_module mux_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
mux_module mux_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
mux_module mux_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
mux_module mux_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
mux_module mux_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
xor_module xor_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
mux_module mux_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
mux_module mux_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
xor_module xor_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
xor_module xor_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
mux_module mux_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
mux_module mux_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
mux_module mux_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
xor_module xor_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
xor_module xor_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
mux_module mux_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
mux_module mux_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
mux_module mux_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
mux_module mux_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [719:0] <= intermediate_reg_1; 
outp[835:720] <= intermediate_reg_1[115:0] ; 
end 
endmodule 
 

module interface_6(input [895:0] inp, output reg [2919:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[895:0] <= inp ; 
outp[1791:896] <= inp ; 
outp[2687:1792] <= inp ; 
outp[2919:2688] <= inp[231:0] ; 
end 
endmodule 

module interface_7(input [2399:0] inp, output reg [3095:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[2399:0] <= inp ; 
outp[3095:2400] <= inp[695:0] ; 
end 
endmodule 

module interface_8(input [2399:0] inp, output reg [3131:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[2399:0] <= inp ; 
outp[3131:2400] <= inp[731:0] ; 
end 
endmodule 

module interface_9(input [1247:0] inp, output reg [895:0] outp, input clk, input reset);
reg [1247:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
wire [623:0]intermediate_reg_1; 
 
xor_module xor_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
xor_module xor_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
xor_module xor_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
xor_module xor_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
xor_module xor_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
mux_module mux_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
xor_module xor_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
xor_module xor_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
xor_module xor_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
mux_module mux_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
xor_module xor_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
xor_module xor_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
mux_module mux_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
xor_module xor_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
mux_module mux_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
xor_module xor_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
mux_module mux_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
mux_module mux_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
mux_module mux_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
mux_module mux_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
mux_module mux_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
xor_module xor_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
mux_module mux_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
xor_module xor_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
mux_module mux_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
mux_module mux_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
mux_module mux_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
mux_module mux_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
mux_module mux_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
mux_module mux_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
mux_module mux_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
mux_module mux_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
xor_module xor_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
xor_module xor_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
xor_module xor_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
xor_module xor_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
mux_module mux_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
xor_module xor_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
xor_module xor_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
xor_module xor_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
mux_module mux_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
xor_module xor_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
xor_module xor_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
xor_module xor_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
xor_module xor_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
xor_module xor_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
mux_module mux_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
xor_module xor_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
xor_module xor_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
mux_module mux_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
xor_module xor_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
mux_module mux_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
xor_module xor_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
xor_module xor_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
xor_module xor_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
xor_module xor_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
mux_module mux_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
mux_module mux_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
xor_module xor_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
mux_module mux_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
xor_module xor_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
xor_module xor_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
xor_module xor_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
xor_module xor_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
xor_module xor_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
mux_module mux_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
xor_module xor_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
xor_module xor_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
mux_module mux_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
xor_module xor_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
xor_module xor_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
mux_module mux_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
mux_module mux_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
mux_module mux_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
xor_module xor_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
mux_module mux_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
xor_module xor_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
mux_module mux_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
mux_module mux_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
xor_module xor_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
xor_module xor_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
mux_module mux_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
mux_module mux_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
mux_module mux_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
xor_module xor_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
mux_module mux_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
mux_module mux_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
mux_module mux_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
xor_module xor_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
xor_module xor_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
mux_module mux_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
xor_module xor_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
mux_module mux_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
xor_module xor_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
mux_module mux_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
xor_module xor_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
mux_module mux_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
xor_module xor_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
mux_module mux_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
xor_module xor_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
xor_module xor_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
xor_module xor_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
xor_module xor_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
xor_module xor_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
xor_module xor_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
xor_module xor_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
mux_module mux_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
mux_module mux_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
mux_module mux_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
xor_module xor_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
xor_module xor_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
xor_module xor_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
mux_module mux_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
xor_module xor_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
xor_module xor_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
mux_module mux_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
mux_module mux_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
mux_module mux_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
mux_module mux_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
mux_module mux_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
xor_module xor_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
xor_module xor_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
mux_module mux_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
xor_module xor_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
xor_module xor_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
mux_module mux_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
xor_module xor_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
xor_module xor_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
mux_module mux_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
xor_module xor_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
xor_module xor_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
xor_module xor_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
xor_module xor_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
xor_module xor_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
xor_module xor_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
mux_module mux_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
xor_module xor_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
xor_module xor_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
xor_module xor_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
xor_module xor_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
xor_module xor_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
xor_module xor_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
mux_module mux_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
mux_module mux_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
xor_module xor_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
xor_module xor_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [623:0] <= intermediate_reg_1; 
outp[895:624] <= intermediate_reg_1[271:0] ; 
end 
endmodule 
 

module interface_10(input [1887:0] inp, output reg [1535:0] outp, input clk, input reset);
reg [1887:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
wire [943:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
xor_module xor_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
mux_module mux_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
mux_module mux_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
xor_module xor_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
xor_module xor_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
xor_module xor_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
xor_module xor_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
xor_module xor_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
xor_module xor_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
xor_module xor_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
xor_module xor_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
mux_module mux_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
xor_module xor_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
xor_module xor_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
xor_module xor_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
mux_module mux_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
xor_module xor_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
mux_module mux_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
mux_module mux_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
mux_module mux_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
xor_module xor_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
xor_module xor_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
mux_module mux_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
mux_module mux_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
xor_module xor_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
xor_module xor_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
xor_module xor_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
xor_module xor_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
xor_module xor_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824])); 
mux_module mux_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
xor_module xor_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810])); 
xor_module xor_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
mux_module mux_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
xor_module xor_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
xor_module xor_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
xor_module xor_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
mux_module mux_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
mux_module mux_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
xor_module xor_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
xor_module xor_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
xor_module xor_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
mux_module mux_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
mux_module mux_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
mux_module mux_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
xor_module xor_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
mux_module mux_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
xor_module xor_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
mux_module mux_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
xor_module xor_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
mux_module mux_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
mux_module mux_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
xor_module xor_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
xor_module xor_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
xor_module xor_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
xor_module xor_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
xor_module xor_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
xor_module xor_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
xor_module xor_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
mux_module mux_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
xor_module xor_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
xor_module xor_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
mux_module mux_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
mux_module mux_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
xor_module xor_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
mux_module mux_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
xor_module xor_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
mux_module mux_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
xor_module xor_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
xor_module xor_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
xor_module xor_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
mux_module mux_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
xor_module xor_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
mux_module mux_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
mux_module mux_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
xor_module xor_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
xor_module xor_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
mux_module mux_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
xor_module xor_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
xor_module xor_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
mux_module mux_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
xor_module xor_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
xor_module xor_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
xor_module xor_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
mux_module mux_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
xor_module xor_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
mux_module mux_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
xor_module xor_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
xor_module xor_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
xor_module xor_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
mux_module mux_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
xor_module xor_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
mux_module mux_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
xor_module xor_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
mux_module mux_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
xor_module xor_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
mux_module mux_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
mux_module mux_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
mux_module mux_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
mux_module mux_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
mux_module mux_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
mux_module mux_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
mux_module mux_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
xor_module xor_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
mux_module mux_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
mux_module mux_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
xor_module xor_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
xor_module xor_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
xor_module xor_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
xor_module xor_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
xor_module xor_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
xor_module xor_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
xor_module xor_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
xor_module xor_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
mux_module mux_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
mux_module mux_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
xor_module xor_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
xor_module xor_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
xor_module xor_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
mux_module mux_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
xor_module xor_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
xor_module xor_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
mux_module mux_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
xor_module xor_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
xor_module xor_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
xor_module xor_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
mux_module mux_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
xor_module xor_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
mux_module mux_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
xor_module xor_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
xor_module xor_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
xor_module xor_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
mux_module mux_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
xor_module xor_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
mux_module mux_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
mux_module mux_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
xor_module xor_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
mux_module mux_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
xor_module xor_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
xor_module xor_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
mux_module mux_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
xor_module xor_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
mux_module mux_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
mux_module mux_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
mux_module mux_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
xor_module xor_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
xor_module xor_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
mux_module mux_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
mux_module mux_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
xor_module xor_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
xor_module xor_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
mux_module mux_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
xor_module xor_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
xor_module xor_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
mux_module mux_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
xor_module xor_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
mux_module mux_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
xor_module xor_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
mux_module mux_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
xor_module xor_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
xor_module xor_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
xor_module xor_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
mux_module mux_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
mux_module mux_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
mux_module mux_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
mux_module mux_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
xor_module xor_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
mux_module mux_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
mux_module mux_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
xor_module xor_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
xor_module xor_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
xor_module xor_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
xor_module xor_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
xor_module xor_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
mux_module mux_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
xor_module xor_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
xor_module xor_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
mux_module mux_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
xor_module xor_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
xor_module xor_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
mux_module mux_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
mux_module mux_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
mux_module mux_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
xor_module xor_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
xor_module xor_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
xor_module xor_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
mux_module mux_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
xor_module xor_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
xor_module xor_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
xor_module xor_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
mux_module mux_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
mux_module mux_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
mux_module mux_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
xor_module xor_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
xor_module xor_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
xor_module xor_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
xor_module xor_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
xor_module xor_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
mux_module mux_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
mux_module mux_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
xor_module xor_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
xor_module xor_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
mux_module mux_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
xor_module xor_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
xor_module xor_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
mux_module mux_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
mux_module mux_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
mux_module mux_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
xor_module xor_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
xor_module xor_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
mux_module mux_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
mux_module mux_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
xor_module xor_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
mux_module mux_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
xor_module xor_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
xor_module xor_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
xor_module xor_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
xor_module xor_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
xor_module xor_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
xor_module xor_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
xor_module xor_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
xor_module xor_module_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
xor_module xor_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
mux_module mux_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
xor_module xor_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
xor_module xor_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
xor_module xor_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
xor_module xor_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
mux_module mux_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
xor_module xor_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
xor_module xor_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
mux_module mux_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
xor_module xor_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
mux_module mux_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
mux_module mux_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
mux_module mux_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
xor_module xor_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
xor_module xor_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
mux_module mux_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
mux_module mux_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
xor_module xor_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
mux_module mux_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
mux_module mux_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
mux_module mux_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
mux_module mux_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
xor_module xor_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
xor_module xor_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
xor_module xor_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
xor_module xor_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
mux_module mux_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
mux_module mux_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
mux_module mux_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
xor_module xor_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
mux_module mux_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
mux_module mux_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
xor_module xor_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
mux_module mux_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
mux_module mux_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
xor_module xor_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
mux_module mux_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
mux_module mux_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
xor_module xor_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
mux_module mux_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
mux_module mux_module_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
xor_module xor_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
mux_module mux_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
mux_module mux_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
xor_module xor_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
mux_module mux_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
xor_module xor_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
xor_module xor_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
mux_module mux_module_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
xor_module xor_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
mux_module mux_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
mux_module mux_module_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
mux_module mux_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
xor_module xor_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
xor_module xor_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
xor_module xor_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
mux_module mux_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
mux_module mux_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
mux_module mux_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
xor_module xor_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
xor_module xor_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
mux_module mux_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
xor_module xor_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
xor_module xor_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
xor_module xor_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
xor_module xor_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
xor_module xor_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
xor_module xor_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
xor_module xor_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
xor_module xor_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
xor_module xor_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
mux_module mux_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
xor_module xor_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
mux_module mux_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
mux_module mux_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
xor_module xor_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
mux_module mux_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
xor_module xor_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
mux_module mux_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
xor_module xor_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
xor_module xor_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
mux_module mux_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
always@(posedge clk) begin 
outp [943:0] <= intermediate_reg_1; 
outp[1535:944] <= intermediate_reg_1[591:0] ; 
end 
endmodule 
 

module interface_11(input [6595:0] inp, output reg [5119:0] outp, input clk, input reset);
reg [6595:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
wire [3297:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6595]),.i2(intermediate_reg_0[6594]),.o(intermediate_reg_1[3297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6593]),.i2(intermediate_reg_0[6592]),.o(intermediate_reg_1[3296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6591]),.i2(intermediate_reg_0[6590]),.o(intermediate_reg_1[3295]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6589]),.i2(intermediate_reg_0[6588]),.o(intermediate_reg_1[3294])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6587]),.i2(intermediate_reg_0[6586]),.o(intermediate_reg_1[3293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6585]),.i2(intermediate_reg_0[6584]),.o(intermediate_reg_1[3292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6583]),.i2(intermediate_reg_0[6582]),.o(intermediate_reg_1[3291]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6581]),.i2(intermediate_reg_0[6580]),.o(intermediate_reg_1[3290]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6579]),.i2(intermediate_reg_0[6578]),.o(intermediate_reg_1[3289])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6577]),.i2(intermediate_reg_0[6576]),.o(intermediate_reg_1[3288]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6575]),.i2(intermediate_reg_0[6574]),.o(intermediate_reg_1[3287])); 
xor_module xor_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6573]),.i2(intermediate_reg_0[6572]),.o(intermediate_reg_1[3286])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6571]),.i2(intermediate_reg_0[6570]),.o(intermediate_reg_1[3285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6569]),.i2(intermediate_reg_0[6568]),.o(intermediate_reg_1[3284]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6567]),.i2(intermediate_reg_0[6566]),.o(intermediate_reg_1[3283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6565]),.i2(intermediate_reg_0[6564]),.o(intermediate_reg_1[3282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6563]),.i2(intermediate_reg_0[6562]),.o(intermediate_reg_1[3281]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6561]),.i2(intermediate_reg_0[6560]),.o(intermediate_reg_1[3280])); 
xor_module xor_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6559]),.i2(intermediate_reg_0[6558]),.o(intermediate_reg_1[3279])); 
xor_module xor_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6557]),.i2(intermediate_reg_0[6556]),.o(intermediate_reg_1[3278])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6555]),.i2(intermediate_reg_0[6554]),.o(intermediate_reg_1[3277])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6553]),.i2(intermediate_reg_0[6552]),.o(intermediate_reg_1[3276]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6551]),.i2(intermediate_reg_0[6550]),.o(intermediate_reg_1[3275])); 
mux_module mux_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6549]),.i2(intermediate_reg_0[6548]),.o(intermediate_reg_1[3274]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6547]),.i2(intermediate_reg_0[6546]),.o(intermediate_reg_1[3273])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6545]),.i2(intermediate_reg_0[6544]),.o(intermediate_reg_1[3272]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6543]),.i2(intermediate_reg_0[6542]),.o(intermediate_reg_1[3271])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6541]),.i2(intermediate_reg_0[6540]),.o(intermediate_reg_1[3270])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6539]),.i2(intermediate_reg_0[6538]),.o(intermediate_reg_1[3269]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6537]),.i2(intermediate_reg_0[6536]),.o(intermediate_reg_1[3268])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6535]),.i2(intermediate_reg_0[6534]),.o(intermediate_reg_1[3267]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6533]),.i2(intermediate_reg_0[6532]),.o(intermediate_reg_1[3266])); 
xor_module xor_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6531]),.i2(intermediate_reg_0[6530]),.o(intermediate_reg_1[3265])); 
mux_module mux_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6529]),.i2(intermediate_reg_0[6528]),.o(intermediate_reg_1[3264]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6527]),.i2(intermediate_reg_0[6526]),.o(intermediate_reg_1[3263]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6525]),.i2(intermediate_reg_0[6524]),.o(intermediate_reg_1[3262])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6523]),.i2(intermediate_reg_0[6522]),.o(intermediate_reg_1[3261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6521]),.i2(intermediate_reg_0[6520]),.o(intermediate_reg_1[3260]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6519]),.i2(intermediate_reg_0[6518]),.o(intermediate_reg_1[3259]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6517]),.i2(intermediate_reg_0[6516]),.o(intermediate_reg_1[3258])); 
mux_module mux_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6515]),.i2(intermediate_reg_0[6514]),.o(intermediate_reg_1[3257]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6513]),.i2(intermediate_reg_0[6512]),.o(intermediate_reg_1[3256]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6511]),.i2(intermediate_reg_0[6510]),.o(intermediate_reg_1[3255])); 
mux_module mux_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6509]),.i2(intermediate_reg_0[6508]),.o(intermediate_reg_1[3254]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6507]),.i2(intermediate_reg_0[6506]),.o(intermediate_reg_1[3253])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6505]),.i2(intermediate_reg_0[6504]),.o(intermediate_reg_1[3252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6503]),.i2(intermediate_reg_0[6502]),.o(intermediate_reg_1[3251]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6501]),.i2(intermediate_reg_0[6500]),.o(intermediate_reg_1[3250]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6499]),.i2(intermediate_reg_0[6498]),.o(intermediate_reg_1[3249]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6497]),.i2(intermediate_reg_0[6496]),.o(intermediate_reg_1[3248])); 
xor_module xor_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6495]),.i2(intermediate_reg_0[6494]),.o(intermediate_reg_1[3247])); 
xor_module xor_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6493]),.i2(intermediate_reg_0[6492]),.o(intermediate_reg_1[3246])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6491]),.i2(intermediate_reg_0[6490]),.o(intermediate_reg_1[3245]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6489]),.i2(intermediate_reg_0[6488]),.o(intermediate_reg_1[3244])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6487]),.i2(intermediate_reg_0[6486]),.o(intermediate_reg_1[3243]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6485]),.i2(intermediate_reg_0[6484]),.o(intermediate_reg_1[3242])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6483]),.i2(intermediate_reg_0[6482]),.o(intermediate_reg_1[3241]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6481]),.i2(intermediate_reg_0[6480]),.o(intermediate_reg_1[3240]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6479]),.i2(intermediate_reg_0[6478]),.o(intermediate_reg_1[3239])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6477]),.i2(intermediate_reg_0[6476]),.o(intermediate_reg_1[3238]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6475]),.i2(intermediate_reg_0[6474]),.o(intermediate_reg_1[3237]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6473]),.i2(intermediate_reg_0[6472]),.o(intermediate_reg_1[3236])); 
xor_module xor_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6471]),.i2(intermediate_reg_0[6470]),.o(intermediate_reg_1[3235])); 
mux_module mux_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6469]),.i2(intermediate_reg_0[6468]),.o(intermediate_reg_1[3234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6467]),.i2(intermediate_reg_0[6466]),.o(intermediate_reg_1[3233]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6465]),.i2(intermediate_reg_0[6464]),.o(intermediate_reg_1[3232])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6463]),.i2(intermediate_reg_0[6462]),.o(intermediate_reg_1[3231]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6461]),.i2(intermediate_reg_0[6460]),.o(intermediate_reg_1[3230])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6459]),.i2(intermediate_reg_0[6458]),.o(intermediate_reg_1[3229]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6457]),.i2(intermediate_reg_0[6456]),.o(intermediate_reg_1[3228])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6455]),.i2(intermediate_reg_0[6454]),.o(intermediate_reg_1[3227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6453]),.i2(intermediate_reg_0[6452]),.o(intermediate_reg_1[3226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6451]),.i2(intermediate_reg_0[6450]),.o(intermediate_reg_1[3225]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6449]),.i2(intermediate_reg_0[6448]),.o(intermediate_reg_1[3224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6447]),.i2(intermediate_reg_0[6446]),.o(intermediate_reg_1[3223]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6445]),.i2(intermediate_reg_0[6444]),.o(intermediate_reg_1[3222]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6443]),.i2(intermediate_reg_0[6442]),.o(intermediate_reg_1[3221])); 
xor_module xor_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6441]),.i2(intermediate_reg_0[6440]),.o(intermediate_reg_1[3220])); 
xor_module xor_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6439]),.i2(intermediate_reg_0[6438]),.o(intermediate_reg_1[3219])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6437]),.i2(intermediate_reg_0[6436]),.o(intermediate_reg_1[3218]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6435]),.i2(intermediate_reg_0[6434]),.o(intermediate_reg_1[3217])); 
mux_module mux_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6433]),.i2(intermediate_reg_0[6432]),.o(intermediate_reg_1[3216]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6431]),.i2(intermediate_reg_0[6430]),.o(intermediate_reg_1[3215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6429]),.i2(intermediate_reg_0[6428]),.o(intermediate_reg_1[3214]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6427]),.i2(intermediate_reg_0[6426]),.o(intermediate_reg_1[3213])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6425]),.i2(intermediate_reg_0[6424]),.o(intermediate_reg_1[3212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6423]),.i2(intermediate_reg_0[6422]),.o(intermediate_reg_1[3211]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6421]),.i2(intermediate_reg_0[6420]),.o(intermediate_reg_1[3210]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6419]),.i2(intermediate_reg_0[6418]),.o(intermediate_reg_1[3209])); 
mux_module mux_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6417]),.i2(intermediate_reg_0[6416]),.o(intermediate_reg_1[3208]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6415]),.i2(intermediate_reg_0[6414]),.o(intermediate_reg_1[3207])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6413]),.i2(intermediate_reg_0[6412]),.o(intermediate_reg_1[3206])); 
mux_module mux_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6411]),.i2(intermediate_reg_0[6410]),.o(intermediate_reg_1[3205]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6409]),.i2(intermediate_reg_0[6408]),.o(intermediate_reg_1[3204])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6407]),.i2(intermediate_reg_0[6406]),.o(intermediate_reg_1[3203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6405]),.i2(intermediate_reg_0[6404]),.o(intermediate_reg_1[3202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6403]),.i2(intermediate_reg_0[6402]),.o(intermediate_reg_1[3201]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6401]),.i2(intermediate_reg_0[6400]),.o(intermediate_reg_1[3200])); 
mux_module mux_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6399]),.i2(intermediate_reg_0[6398]),.o(intermediate_reg_1[3199]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6397]),.i2(intermediate_reg_0[6396]),.o(intermediate_reg_1[3198]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6395]),.i2(intermediate_reg_0[6394]),.o(intermediate_reg_1[3197])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6393]),.i2(intermediate_reg_0[6392]),.o(intermediate_reg_1[3196])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6391]),.i2(intermediate_reg_0[6390]),.o(intermediate_reg_1[3195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6389]),.i2(intermediate_reg_0[6388]),.o(intermediate_reg_1[3194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6387]),.i2(intermediate_reg_0[6386]),.o(intermediate_reg_1[3193]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6385]),.i2(intermediate_reg_0[6384]),.o(intermediate_reg_1[3192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6383]),.i2(intermediate_reg_0[6382]),.o(intermediate_reg_1[3191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6381]),.i2(intermediate_reg_0[6380]),.o(intermediate_reg_1[3190]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6379]),.i2(intermediate_reg_0[6378]),.o(intermediate_reg_1[3189])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6377]),.i2(intermediate_reg_0[6376]),.o(intermediate_reg_1[3188])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6375]),.i2(intermediate_reg_0[6374]),.o(intermediate_reg_1[3187])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6373]),.i2(intermediate_reg_0[6372]),.o(intermediate_reg_1[3186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6371]),.i2(intermediate_reg_0[6370]),.o(intermediate_reg_1[3185]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6369]),.i2(intermediate_reg_0[6368]),.o(intermediate_reg_1[3184])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6367]),.i2(intermediate_reg_0[6366]),.o(intermediate_reg_1[3183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6365]),.i2(intermediate_reg_0[6364]),.o(intermediate_reg_1[3182]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6363]),.i2(intermediate_reg_0[6362]),.o(intermediate_reg_1[3181]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6361]),.i2(intermediate_reg_0[6360]),.o(intermediate_reg_1[3180])); 
mux_module mux_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6359]),.i2(intermediate_reg_0[6358]),.o(intermediate_reg_1[3179]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6357]),.i2(intermediate_reg_0[6356]),.o(intermediate_reg_1[3178])); 
mux_module mux_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6355]),.i2(intermediate_reg_0[6354]),.o(intermediate_reg_1[3177]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6353]),.i2(intermediate_reg_0[6352]),.o(intermediate_reg_1[3176])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6351]),.i2(intermediate_reg_0[6350]),.o(intermediate_reg_1[3175]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6349]),.i2(intermediate_reg_0[6348]),.o(intermediate_reg_1[3174])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6347]),.i2(intermediate_reg_0[6346]),.o(intermediate_reg_1[3173])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6345]),.i2(intermediate_reg_0[6344]),.o(intermediate_reg_1[3172])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6343]),.i2(intermediate_reg_0[6342]),.o(intermediate_reg_1[3171]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6341]),.i2(intermediate_reg_0[6340]),.o(intermediate_reg_1[3170])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6339]),.i2(intermediate_reg_0[6338]),.o(intermediate_reg_1[3169]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6337]),.i2(intermediate_reg_0[6336]),.o(intermediate_reg_1[3168])); 
mux_module mux_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6335]),.i2(intermediate_reg_0[6334]),.o(intermediate_reg_1[3167]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6333]),.i2(intermediate_reg_0[6332]),.o(intermediate_reg_1[3166])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6331]),.i2(intermediate_reg_0[6330]),.o(intermediate_reg_1[3165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6329]),.i2(intermediate_reg_0[6328]),.o(intermediate_reg_1[3164])); 
xor_module xor_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6327]),.i2(intermediate_reg_0[6326]),.o(intermediate_reg_1[3163])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6325]),.i2(intermediate_reg_0[6324]),.o(intermediate_reg_1[3162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6323]),.i2(intermediate_reg_0[6322]),.o(intermediate_reg_1[3161]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6321]),.i2(intermediate_reg_0[6320]),.o(intermediate_reg_1[3160])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6319]),.i2(intermediate_reg_0[6318]),.o(intermediate_reg_1[3159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6317]),.i2(intermediate_reg_0[6316]),.o(intermediate_reg_1[3158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6315]),.i2(intermediate_reg_0[6314]),.o(intermediate_reg_1[3157]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6313]),.i2(intermediate_reg_0[6312]),.o(intermediate_reg_1[3156])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6311]),.i2(intermediate_reg_0[6310]),.o(intermediate_reg_1[3155])); 
xor_module xor_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6309]),.i2(intermediate_reg_0[6308]),.o(intermediate_reg_1[3154])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6307]),.i2(intermediate_reg_0[6306]),.o(intermediate_reg_1[3153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6305]),.i2(intermediate_reg_0[6304]),.o(intermediate_reg_1[3152]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6303]),.i2(intermediate_reg_0[6302]),.o(intermediate_reg_1[3151])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6301]),.i2(intermediate_reg_0[6300]),.o(intermediate_reg_1[3150])); 
xor_module xor_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6299]),.i2(intermediate_reg_0[6298]),.o(intermediate_reg_1[3149])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6297]),.i2(intermediate_reg_0[6296]),.o(intermediate_reg_1[3148]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6295]),.i2(intermediate_reg_0[6294]),.o(intermediate_reg_1[3147])); 
xor_module xor_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6293]),.i2(intermediate_reg_0[6292]),.o(intermediate_reg_1[3146])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6291]),.i2(intermediate_reg_0[6290]),.o(intermediate_reg_1[3145])); 
xor_module xor_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6289]),.i2(intermediate_reg_0[6288]),.o(intermediate_reg_1[3144])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6287]),.i2(intermediate_reg_0[6286]),.o(intermediate_reg_1[3143]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6285]),.i2(intermediate_reg_0[6284]),.o(intermediate_reg_1[3142])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6283]),.i2(intermediate_reg_0[6282]),.o(intermediate_reg_1[3141]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6281]),.i2(intermediate_reg_0[6280]),.o(intermediate_reg_1[3140])); 
mux_module mux_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6279]),.i2(intermediate_reg_0[6278]),.o(intermediate_reg_1[3139]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6277]),.i2(intermediate_reg_0[6276]),.o(intermediate_reg_1[3138])); 
mux_module mux_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6275]),.i2(intermediate_reg_0[6274]),.o(intermediate_reg_1[3137]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6273]),.i2(intermediate_reg_0[6272]),.o(intermediate_reg_1[3136]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6271]),.i2(intermediate_reg_0[6270]),.o(intermediate_reg_1[3135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6269]),.i2(intermediate_reg_0[6268]),.o(intermediate_reg_1[3134]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6267]),.i2(intermediate_reg_0[6266]),.o(intermediate_reg_1[3133])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6265]),.i2(intermediate_reg_0[6264]),.o(intermediate_reg_1[3132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6263]),.i2(intermediate_reg_0[6262]),.o(intermediate_reg_1[3131]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6261]),.i2(intermediate_reg_0[6260]),.o(intermediate_reg_1[3130])); 
xor_module xor_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6259]),.i2(intermediate_reg_0[6258]),.o(intermediate_reg_1[3129])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6257]),.i2(intermediate_reg_0[6256]),.o(intermediate_reg_1[3128])); 
xor_module xor_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6255]),.i2(intermediate_reg_0[6254]),.o(intermediate_reg_1[3127])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6253]),.i2(intermediate_reg_0[6252]),.o(intermediate_reg_1[3126]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6251]),.i2(intermediate_reg_0[6250]),.o(intermediate_reg_1[3125]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6249]),.i2(intermediate_reg_0[6248]),.o(intermediate_reg_1[3124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6247]),.i2(intermediate_reg_0[6246]),.o(intermediate_reg_1[3123]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6245]),.i2(intermediate_reg_0[6244]),.o(intermediate_reg_1[3122])); 
xor_module xor_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6243]),.i2(intermediate_reg_0[6242]),.o(intermediate_reg_1[3121])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6241]),.i2(intermediate_reg_0[6240]),.o(intermediate_reg_1[3120])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6239]),.i2(intermediate_reg_0[6238]),.o(intermediate_reg_1[3119])); 
xor_module xor_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6237]),.i2(intermediate_reg_0[6236]),.o(intermediate_reg_1[3118])); 
mux_module mux_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6235]),.i2(intermediate_reg_0[6234]),.o(intermediate_reg_1[3117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6233]),.i2(intermediate_reg_0[6232]),.o(intermediate_reg_1[3116]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6231]),.i2(intermediate_reg_0[6230]),.o(intermediate_reg_1[3115])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6229]),.i2(intermediate_reg_0[6228]),.o(intermediate_reg_1[3114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6227]),.i2(intermediate_reg_0[6226]),.o(intermediate_reg_1[3113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6225]),.i2(intermediate_reg_0[6224]),.o(intermediate_reg_1[3112]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6223]),.i2(intermediate_reg_0[6222]),.o(intermediate_reg_1[3111])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6221]),.i2(intermediate_reg_0[6220]),.o(intermediate_reg_1[3110]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6219]),.i2(intermediate_reg_0[6218]),.o(intermediate_reg_1[3109])); 
xor_module xor_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6217]),.i2(intermediate_reg_0[6216]),.o(intermediate_reg_1[3108])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6215]),.i2(intermediate_reg_0[6214]),.o(intermediate_reg_1[3107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6213]),.i2(intermediate_reg_0[6212]),.o(intermediate_reg_1[3106]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6211]),.i2(intermediate_reg_0[6210]),.o(intermediate_reg_1[3105]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6209]),.i2(intermediate_reg_0[6208]),.o(intermediate_reg_1[3104])); 
xor_module xor_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6207]),.i2(intermediate_reg_0[6206]),.o(intermediate_reg_1[3103])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6205]),.i2(intermediate_reg_0[6204]),.o(intermediate_reg_1[3102]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6203]),.i2(intermediate_reg_0[6202]),.o(intermediate_reg_1[3101])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6201]),.i2(intermediate_reg_0[6200]),.o(intermediate_reg_1[3100]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6199]),.i2(intermediate_reg_0[6198]),.o(intermediate_reg_1[3099])); 
xor_module xor_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6197]),.i2(intermediate_reg_0[6196]),.o(intermediate_reg_1[3098])); 
xor_module xor_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6195]),.i2(intermediate_reg_0[6194]),.o(intermediate_reg_1[3097])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6193]),.i2(intermediate_reg_0[6192]),.o(intermediate_reg_1[3096]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6191]),.i2(intermediate_reg_0[6190]),.o(intermediate_reg_1[3095]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6189]),.i2(intermediate_reg_0[6188]),.o(intermediate_reg_1[3094]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6187]),.i2(intermediate_reg_0[6186]),.o(intermediate_reg_1[3093])); 
xor_module xor_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6185]),.i2(intermediate_reg_0[6184]),.o(intermediate_reg_1[3092])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6183]),.i2(intermediate_reg_0[6182]),.o(intermediate_reg_1[3091]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6181]),.i2(intermediate_reg_0[6180]),.o(intermediate_reg_1[3090]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6179]),.i2(intermediate_reg_0[6178]),.o(intermediate_reg_1[3089]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6177]),.i2(intermediate_reg_0[6176]),.o(intermediate_reg_1[3088])); 
mux_module mux_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6175]),.i2(intermediate_reg_0[6174]),.o(intermediate_reg_1[3087]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6173]),.i2(intermediate_reg_0[6172]),.o(intermediate_reg_1[3086])); 
xor_module xor_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6171]),.i2(intermediate_reg_0[6170]),.o(intermediate_reg_1[3085])); 
xor_module xor_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6169]),.i2(intermediate_reg_0[6168]),.o(intermediate_reg_1[3084])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6167]),.i2(intermediate_reg_0[6166]),.o(intermediate_reg_1[3083]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6165]),.i2(intermediate_reg_0[6164]),.o(intermediate_reg_1[3082])); 
mux_module mux_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6163]),.i2(intermediate_reg_0[6162]),.o(intermediate_reg_1[3081]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6161]),.i2(intermediate_reg_0[6160]),.o(intermediate_reg_1[3080]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6159]),.i2(intermediate_reg_0[6158]),.o(intermediate_reg_1[3079]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6157]),.i2(intermediate_reg_0[6156]),.o(intermediate_reg_1[3078]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6155]),.i2(intermediate_reg_0[6154]),.o(intermediate_reg_1[3077])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6153]),.i2(intermediate_reg_0[6152]),.o(intermediate_reg_1[3076]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6151]),.i2(intermediate_reg_0[6150]),.o(intermediate_reg_1[3075]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6149]),.i2(intermediate_reg_0[6148]),.o(intermediate_reg_1[3074]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6147]),.i2(intermediate_reg_0[6146]),.o(intermediate_reg_1[3073])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6145]),.i2(intermediate_reg_0[6144]),.o(intermediate_reg_1[3072]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6143]),.i2(intermediate_reg_0[6142]),.o(intermediate_reg_1[3071])); 
mux_module mux_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6141]),.i2(intermediate_reg_0[6140]),.o(intermediate_reg_1[3070]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6139]),.i2(intermediate_reg_0[6138]),.o(intermediate_reg_1[3069]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6137]),.i2(intermediate_reg_0[6136]),.o(intermediate_reg_1[3068]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6135]),.i2(intermediate_reg_0[6134]),.o(intermediate_reg_1[3067])); 
xor_module xor_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6133]),.i2(intermediate_reg_0[6132]),.o(intermediate_reg_1[3066])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6131]),.i2(intermediate_reg_0[6130]),.o(intermediate_reg_1[3065])); 
xor_module xor_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6129]),.i2(intermediate_reg_0[6128]),.o(intermediate_reg_1[3064])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6127]),.i2(intermediate_reg_0[6126]),.o(intermediate_reg_1[3063])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6125]),.i2(intermediate_reg_0[6124]),.o(intermediate_reg_1[3062]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6123]),.i2(intermediate_reg_0[6122]),.o(intermediate_reg_1[3061])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6121]),.i2(intermediate_reg_0[6120]),.o(intermediate_reg_1[3060])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6119]),.i2(intermediate_reg_0[6118]),.o(intermediate_reg_1[3059]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6117]),.i2(intermediate_reg_0[6116]),.o(intermediate_reg_1[3058])); 
xor_module xor_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6115]),.i2(intermediate_reg_0[6114]),.o(intermediate_reg_1[3057])); 
mux_module mux_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6113]),.i2(intermediate_reg_0[6112]),.o(intermediate_reg_1[3056]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6111]),.i2(intermediate_reg_0[6110]),.o(intermediate_reg_1[3055])); 
mux_module mux_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6109]),.i2(intermediate_reg_0[6108]),.o(intermediate_reg_1[3054]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6107]),.i2(intermediate_reg_0[6106]),.o(intermediate_reg_1[3053])); 
xor_module xor_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6105]),.i2(intermediate_reg_0[6104]),.o(intermediate_reg_1[3052])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6103]),.i2(intermediate_reg_0[6102]),.o(intermediate_reg_1[3051]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6101]),.i2(intermediate_reg_0[6100]),.o(intermediate_reg_1[3050]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6099]),.i2(intermediate_reg_0[6098]),.o(intermediate_reg_1[3049])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6097]),.i2(intermediate_reg_0[6096]),.o(intermediate_reg_1[3048]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6095]),.i2(intermediate_reg_0[6094]),.o(intermediate_reg_1[3047]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6093]),.i2(intermediate_reg_0[6092]),.o(intermediate_reg_1[3046]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6091]),.i2(intermediate_reg_0[6090]),.o(intermediate_reg_1[3045])); 
xor_module xor_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6089]),.i2(intermediate_reg_0[6088]),.o(intermediate_reg_1[3044])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6087]),.i2(intermediate_reg_0[6086]),.o(intermediate_reg_1[3043]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6085]),.i2(intermediate_reg_0[6084]),.o(intermediate_reg_1[3042]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6083]),.i2(intermediate_reg_0[6082]),.o(intermediate_reg_1[3041]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6081]),.i2(intermediate_reg_0[6080]),.o(intermediate_reg_1[3040]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6079]),.i2(intermediate_reg_0[6078]),.o(intermediate_reg_1[3039]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6077]),.i2(intermediate_reg_0[6076]),.o(intermediate_reg_1[3038]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6075]),.i2(intermediate_reg_0[6074]),.o(intermediate_reg_1[3037])); 
xor_module xor_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6073]),.i2(intermediate_reg_0[6072]),.o(intermediate_reg_1[3036])); 
xor_module xor_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6071]),.i2(intermediate_reg_0[6070]),.o(intermediate_reg_1[3035])); 
xor_module xor_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6069]),.i2(intermediate_reg_0[6068]),.o(intermediate_reg_1[3034])); 
xor_module xor_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6067]),.i2(intermediate_reg_0[6066]),.o(intermediate_reg_1[3033])); 
xor_module xor_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6065]),.i2(intermediate_reg_0[6064]),.o(intermediate_reg_1[3032])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6063]),.i2(intermediate_reg_0[6062]),.o(intermediate_reg_1[3031]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6061]),.i2(intermediate_reg_0[6060]),.o(intermediate_reg_1[3030]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6059]),.i2(intermediate_reg_0[6058]),.o(intermediate_reg_1[3029])); 
mux_module mux_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6057]),.i2(intermediate_reg_0[6056]),.o(intermediate_reg_1[3028]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6055]),.i2(intermediate_reg_0[6054]),.o(intermediate_reg_1[3027])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6053]),.i2(intermediate_reg_0[6052]),.o(intermediate_reg_1[3026])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6051]),.i2(intermediate_reg_0[6050]),.o(intermediate_reg_1[3025]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6049]),.i2(intermediate_reg_0[6048]),.o(intermediate_reg_1[3024])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6047]),.i2(intermediate_reg_0[6046]),.o(intermediate_reg_1[3023]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6045]),.i2(intermediate_reg_0[6044]),.o(intermediate_reg_1[3022])); 
xor_module xor_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6043]),.i2(intermediate_reg_0[6042]),.o(intermediate_reg_1[3021])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6041]),.i2(intermediate_reg_0[6040]),.o(intermediate_reg_1[3020])); 
xor_module xor_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6039]),.i2(intermediate_reg_0[6038]),.o(intermediate_reg_1[3019])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6037]),.i2(intermediate_reg_0[6036]),.o(intermediate_reg_1[3018]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6035]),.i2(intermediate_reg_0[6034]),.o(intermediate_reg_1[3017])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6033]),.i2(intermediate_reg_0[6032]),.o(intermediate_reg_1[3016]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6031]),.i2(intermediate_reg_0[6030]),.o(intermediate_reg_1[3015])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6029]),.i2(intermediate_reg_0[6028]),.o(intermediate_reg_1[3014])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6027]),.i2(intermediate_reg_0[6026]),.o(intermediate_reg_1[3013]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6025]),.i2(intermediate_reg_0[6024]),.o(intermediate_reg_1[3012]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6023]),.i2(intermediate_reg_0[6022]),.o(intermediate_reg_1[3011])); 
mux_module mux_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6021]),.i2(intermediate_reg_0[6020]),.o(intermediate_reg_1[3010]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6019]),.i2(intermediate_reg_0[6018]),.o(intermediate_reg_1[3009])); 
xor_module xor_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6017]),.i2(intermediate_reg_0[6016]),.o(intermediate_reg_1[3008])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6015]),.i2(intermediate_reg_0[6014]),.o(intermediate_reg_1[3007])); 
xor_module xor_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6013]),.i2(intermediate_reg_0[6012]),.o(intermediate_reg_1[3006])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6011]),.i2(intermediate_reg_0[6010]),.o(intermediate_reg_1[3005]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6009]),.i2(intermediate_reg_0[6008]),.o(intermediate_reg_1[3004])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6007]),.i2(intermediate_reg_0[6006]),.o(intermediate_reg_1[3003]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6005]),.i2(intermediate_reg_0[6004]),.o(intermediate_reg_1[3002]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6003]),.i2(intermediate_reg_0[6002]),.o(intermediate_reg_1[3001]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6001]),.i2(intermediate_reg_0[6000]),.o(intermediate_reg_1[3000]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5999]),.i2(intermediate_reg_0[5998]),.o(intermediate_reg_1[2999])); 
mux_module mux_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5997]),.i2(intermediate_reg_0[5996]),.o(intermediate_reg_1[2998]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5995]),.i2(intermediate_reg_0[5994]),.o(intermediate_reg_1[2997])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5993]),.i2(intermediate_reg_0[5992]),.o(intermediate_reg_1[2996]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5991]),.i2(intermediate_reg_0[5990]),.o(intermediate_reg_1[2995])); 
mux_module mux_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5989]),.i2(intermediate_reg_0[5988]),.o(intermediate_reg_1[2994]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5987]),.i2(intermediate_reg_0[5986]),.o(intermediate_reg_1[2993]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5985]),.i2(intermediate_reg_0[5984]),.o(intermediate_reg_1[2992])); 
mux_module mux_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5983]),.i2(intermediate_reg_0[5982]),.o(intermediate_reg_1[2991]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5981]),.i2(intermediate_reg_0[5980]),.o(intermediate_reg_1[2990])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5979]),.i2(intermediate_reg_0[5978]),.o(intermediate_reg_1[2989])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5977]),.i2(intermediate_reg_0[5976]),.o(intermediate_reg_1[2988]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5975]),.i2(intermediate_reg_0[5974]),.o(intermediate_reg_1[2987]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5973]),.i2(intermediate_reg_0[5972]),.o(intermediate_reg_1[2986])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5971]),.i2(intermediate_reg_0[5970]),.o(intermediate_reg_1[2985])); 
mux_module mux_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5969]),.i2(intermediate_reg_0[5968]),.o(intermediate_reg_1[2984]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5967]),.i2(intermediate_reg_0[5966]),.o(intermediate_reg_1[2983])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5965]),.i2(intermediate_reg_0[5964]),.o(intermediate_reg_1[2982])); 
mux_module mux_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5963]),.i2(intermediate_reg_0[5962]),.o(intermediate_reg_1[2981]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5961]),.i2(intermediate_reg_0[5960]),.o(intermediate_reg_1[2980])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5959]),.i2(intermediate_reg_0[5958]),.o(intermediate_reg_1[2979])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5957]),.i2(intermediate_reg_0[5956]),.o(intermediate_reg_1[2978])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5955]),.i2(intermediate_reg_0[5954]),.o(intermediate_reg_1[2977]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5953]),.i2(intermediate_reg_0[5952]),.o(intermediate_reg_1[2976]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5951]),.i2(intermediate_reg_0[5950]),.o(intermediate_reg_1[2975])); 
xor_module xor_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5949]),.i2(intermediate_reg_0[5948]),.o(intermediate_reg_1[2974])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5947]),.i2(intermediate_reg_0[5946]),.o(intermediate_reg_1[2973])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5945]),.i2(intermediate_reg_0[5944]),.o(intermediate_reg_1[2972])); 
xor_module xor_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5943]),.i2(intermediate_reg_0[5942]),.o(intermediate_reg_1[2971])); 
xor_module xor_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5941]),.i2(intermediate_reg_0[5940]),.o(intermediate_reg_1[2970])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5939]),.i2(intermediate_reg_0[5938]),.o(intermediate_reg_1[2969])); 
mux_module mux_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5937]),.i2(intermediate_reg_0[5936]),.o(intermediate_reg_1[2968]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5935]),.i2(intermediate_reg_0[5934]),.o(intermediate_reg_1[2967]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5933]),.i2(intermediate_reg_0[5932]),.o(intermediate_reg_1[2966]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5931]),.i2(intermediate_reg_0[5930]),.o(intermediate_reg_1[2965]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5929]),.i2(intermediate_reg_0[5928]),.o(intermediate_reg_1[2964]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5927]),.i2(intermediate_reg_0[5926]),.o(intermediate_reg_1[2963]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5925]),.i2(intermediate_reg_0[5924]),.o(intermediate_reg_1[2962])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5923]),.i2(intermediate_reg_0[5922]),.o(intermediate_reg_1[2961])); 
xor_module xor_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5921]),.i2(intermediate_reg_0[5920]),.o(intermediate_reg_1[2960])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5919]),.i2(intermediate_reg_0[5918]),.o(intermediate_reg_1[2959])); 
mux_module mux_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5917]),.i2(intermediate_reg_0[5916]),.o(intermediate_reg_1[2958]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5915]),.i2(intermediate_reg_0[5914]),.o(intermediate_reg_1[2957])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5913]),.i2(intermediate_reg_0[5912]),.o(intermediate_reg_1[2956])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5911]),.i2(intermediate_reg_0[5910]),.o(intermediate_reg_1[2955]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5909]),.i2(intermediate_reg_0[5908]),.o(intermediate_reg_1[2954]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5907]),.i2(intermediate_reg_0[5906]),.o(intermediate_reg_1[2953]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5905]),.i2(intermediate_reg_0[5904]),.o(intermediate_reg_1[2952])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5903]),.i2(intermediate_reg_0[5902]),.o(intermediate_reg_1[2951])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5901]),.i2(intermediate_reg_0[5900]),.o(intermediate_reg_1[2950])); 
xor_module xor_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5899]),.i2(intermediate_reg_0[5898]),.o(intermediate_reg_1[2949])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5897]),.i2(intermediate_reg_0[5896]),.o(intermediate_reg_1[2948]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5895]),.i2(intermediate_reg_0[5894]),.o(intermediate_reg_1[2947])); 
xor_module xor_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5893]),.i2(intermediate_reg_0[5892]),.o(intermediate_reg_1[2946])); 
xor_module xor_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5891]),.i2(intermediate_reg_0[5890]),.o(intermediate_reg_1[2945])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5889]),.i2(intermediate_reg_0[5888]),.o(intermediate_reg_1[2944])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5887]),.i2(intermediate_reg_0[5886]),.o(intermediate_reg_1[2943])); 
xor_module xor_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5885]),.i2(intermediate_reg_0[5884]),.o(intermediate_reg_1[2942])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5883]),.i2(intermediate_reg_0[5882]),.o(intermediate_reg_1[2941])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5881]),.i2(intermediate_reg_0[5880]),.o(intermediate_reg_1[2940]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5879]),.i2(intermediate_reg_0[5878]),.o(intermediate_reg_1[2939]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5877]),.i2(intermediate_reg_0[5876]),.o(intermediate_reg_1[2938]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5875]),.i2(intermediate_reg_0[5874]),.o(intermediate_reg_1[2937])); 
mux_module mux_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5873]),.i2(intermediate_reg_0[5872]),.o(intermediate_reg_1[2936]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5871]),.i2(intermediate_reg_0[5870]),.o(intermediate_reg_1[2935])); 
mux_module mux_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5869]),.i2(intermediate_reg_0[5868]),.o(intermediate_reg_1[2934]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5867]),.i2(intermediate_reg_0[5866]),.o(intermediate_reg_1[2933])); 
xor_module xor_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5865]),.i2(intermediate_reg_0[5864]),.o(intermediate_reg_1[2932])); 
mux_module mux_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5863]),.i2(intermediate_reg_0[5862]),.o(intermediate_reg_1[2931]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5861]),.i2(intermediate_reg_0[5860]),.o(intermediate_reg_1[2930])); 
xor_module xor_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5859]),.i2(intermediate_reg_0[5858]),.o(intermediate_reg_1[2929])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5857]),.i2(intermediate_reg_0[5856]),.o(intermediate_reg_1[2928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5855]),.i2(intermediate_reg_0[5854]),.o(intermediate_reg_1[2927]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5853]),.i2(intermediate_reg_0[5852]),.o(intermediate_reg_1[2926])); 
mux_module mux_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5851]),.i2(intermediate_reg_0[5850]),.o(intermediate_reg_1[2925]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5849]),.i2(intermediate_reg_0[5848]),.o(intermediate_reg_1[2924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5847]),.i2(intermediate_reg_0[5846]),.o(intermediate_reg_1[2923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5845]),.i2(intermediate_reg_0[5844]),.o(intermediate_reg_1[2922]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5843]),.i2(intermediate_reg_0[5842]),.o(intermediate_reg_1[2921])); 
xor_module xor_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5841]),.i2(intermediate_reg_0[5840]),.o(intermediate_reg_1[2920])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5839]),.i2(intermediate_reg_0[5838]),.o(intermediate_reg_1[2919])); 
mux_module mux_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5837]),.i2(intermediate_reg_0[5836]),.o(intermediate_reg_1[2918]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5835]),.i2(intermediate_reg_0[5834]),.o(intermediate_reg_1[2917]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5833]),.i2(intermediate_reg_0[5832]),.o(intermediate_reg_1[2916]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5831]),.i2(intermediate_reg_0[5830]),.o(intermediate_reg_1[2915]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5829]),.i2(intermediate_reg_0[5828]),.o(intermediate_reg_1[2914]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5827]),.i2(intermediate_reg_0[5826]),.o(intermediate_reg_1[2913])); 
xor_module xor_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5825]),.i2(intermediate_reg_0[5824]),.o(intermediate_reg_1[2912])); 
xor_module xor_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5823]),.i2(intermediate_reg_0[5822]),.o(intermediate_reg_1[2911])); 
xor_module xor_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5821]),.i2(intermediate_reg_0[5820]),.o(intermediate_reg_1[2910])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5819]),.i2(intermediate_reg_0[5818]),.o(intermediate_reg_1[2909])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5817]),.i2(intermediate_reg_0[5816]),.o(intermediate_reg_1[2908]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5815]),.i2(intermediate_reg_0[5814]),.o(intermediate_reg_1[2907]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5813]),.i2(intermediate_reg_0[5812]),.o(intermediate_reg_1[2906])); 
xor_module xor_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5811]),.i2(intermediate_reg_0[5810]),.o(intermediate_reg_1[2905])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5809]),.i2(intermediate_reg_0[5808]),.o(intermediate_reg_1[2904]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5807]),.i2(intermediate_reg_0[5806]),.o(intermediate_reg_1[2903]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5805]),.i2(intermediate_reg_0[5804]),.o(intermediate_reg_1[2902])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5803]),.i2(intermediate_reg_0[5802]),.o(intermediate_reg_1[2901]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5801]),.i2(intermediate_reg_0[5800]),.o(intermediate_reg_1[2900]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5799]),.i2(intermediate_reg_0[5798]),.o(intermediate_reg_1[2899])); 
mux_module mux_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5797]),.i2(intermediate_reg_0[5796]),.o(intermediate_reg_1[2898]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5795]),.i2(intermediate_reg_0[5794]),.o(intermediate_reg_1[2897])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5793]),.i2(intermediate_reg_0[5792]),.o(intermediate_reg_1[2896]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5791]),.i2(intermediate_reg_0[5790]),.o(intermediate_reg_1[2895])); 
mux_module mux_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5789]),.i2(intermediate_reg_0[5788]),.o(intermediate_reg_1[2894]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5787]),.i2(intermediate_reg_0[5786]),.o(intermediate_reg_1[2893])); 
mux_module mux_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5785]),.i2(intermediate_reg_0[5784]),.o(intermediate_reg_1[2892]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5783]),.i2(intermediate_reg_0[5782]),.o(intermediate_reg_1[2891])); 
mux_module mux_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5781]),.i2(intermediate_reg_0[5780]),.o(intermediate_reg_1[2890]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5779]),.i2(intermediate_reg_0[5778]),.o(intermediate_reg_1[2889]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5777]),.i2(intermediate_reg_0[5776]),.o(intermediate_reg_1[2888])); 
xor_module xor_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5775]),.i2(intermediate_reg_0[5774]),.o(intermediate_reg_1[2887])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5773]),.i2(intermediate_reg_0[5772]),.o(intermediate_reg_1[2886])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5771]),.i2(intermediate_reg_0[5770]),.o(intermediate_reg_1[2885])); 
xor_module xor_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5769]),.i2(intermediate_reg_0[5768]),.o(intermediate_reg_1[2884])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5767]),.i2(intermediate_reg_0[5766]),.o(intermediate_reg_1[2883]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5765]),.i2(intermediate_reg_0[5764]),.o(intermediate_reg_1[2882])); 
mux_module mux_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5763]),.i2(intermediate_reg_0[5762]),.o(intermediate_reg_1[2881]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5761]),.i2(intermediate_reg_0[5760]),.o(intermediate_reg_1[2880]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5759]),.i2(intermediate_reg_0[5758]),.o(intermediate_reg_1[2879])); 
mux_module mux_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5757]),.i2(intermediate_reg_0[5756]),.o(intermediate_reg_1[2878]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5755]),.i2(intermediate_reg_0[5754]),.o(intermediate_reg_1[2877])); 
mux_module mux_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5753]),.i2(intermediate_reg_0[5752]),.o(intermediate_reg_1[2876]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5751]),.i2(intermediate_reg_0[5750]),.o(intermediate_reg_1[2875])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5749]),.i2(intermediate_reg_0[5748]),.o(intermediate_reg_1[2874]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5747]),.i2(intermediate_reg_0[5746]),.o(intermediate_reg_1[2873])); 
mux_module mux_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5745]),.i2(intermediate_reg_0[5744]),.o(intermediate_reg_1[2872]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5743]),.i2(intermediate_reg_0[5742]),.o(intermediate_reg_1[2871])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5741]),.i2(intermediate_reg_0[5740]),.o(intermediate_reg_1[2870]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5739]),.i2(intermediate_reg_0[5738]),.o(intermediate_reg_1[2869]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5737]),.i2(intermediate_reg_0[5736]),.o(intermediate_reg_1[2868]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5735]),.i2(intermediate_reg_0[5734]),.o(intermediate_reg_1[2867])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5733]),.i2(intermediate_reg_0[5732]),.o(intermediate_reg_1[2866]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5731]),.i2(intermediate_reg_0[5730]),.o(intermediate_reg_1[2865]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5729]),.i2(intermediate_reg_0[5728]),.o(intermediate_reg_1[2864])); 
xor_module xor_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5727]),.i2(intermediate_reg_0[5726]),.o(intermediate_reg_1[2863])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5725]),.i2(intermediate_reg_0[5724]),.o(intermediate_reg_1[2862])); 
xor_module xor_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5723]),.i2(intermediate_reg_0[5722]),.o(intermediate_reg_1[2861])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5721]),.i2(intermediate_reg_0[5720]),.o(intermediate_reg_1[2860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5719]),.i2(intermediate_reg_0[5718]),.o(intermediate_reg_1[2859]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5717]),.i2(intermediate_reg_0[5716]),.o(intermediate_reg_1[2858])); 
xor_module xor_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5715]),.i2(intermediate_reg_0[5714]),.o(intermediate_reg_1[2857])); 
mux_module mux_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5713]),.i2(intermediate_reg_0[5712]),.o(intermediate_reg_1[2856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5711]),.i2(intermediate_reg_0[5710]),.o(intermediate_reg_1[2855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5709]),.i2(intermediate_reg_0[5708]),.o(intermediate_reg_1[2854]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5707]),.i2(intermediate_reg_0[5706]),.o(intermediate_reg_1[2853])); 
mux_module mux_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5705]),.i2(intermediate_reg_0[5704]),.o(intermediate_reg_1[2852]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5703]),.i2(intermediate_reg_0[5702]),.o(intermediate_reg_1[2851])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5701]),.i2(intermediate_reg_0[5700]),.o(intermediate_reg_1[2850])); 
mux_module mux_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5699]),.i2(intermediate_reg_0[5698]),.o(intermediate_reg_1[2849]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5697]),.i2(intermediate_reg_0[5696]),.o(intermediate_reg_1[2848]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5695]),.i2(intermediate_reg_0[5694]),.o(intermediate_reg_1[2847]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5693]),.i2(intermediate_reg_0[5692]),.o(intermediate_reg_1[2846]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5691]),.i2(intermediate_reg_0[5690]),.o(intermediate_reg_1[2845]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5689]),.i2(intermediate_reg_0[5688]),.o(intermediate_reg_1[2844]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5687]),.i2(intermediate_reg_0[5686]),.o(intermediate_reg_1[2843]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5685]),.i2(intermediate_reg_0[5684]),.o(intermediate_reg_1[2842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5683]),.i2(intermediate_reg_0[5682]),.o(intermediate_reg_1[2841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5681]),.i2(intermediate_reg_0[5680]),.o(intermediate_reg_1[2840]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5679]),.i2(intermediate_reg_0[5678]),.o(intermediate_reg_1[2839])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5677]),.i2(intermediate_reg_0[5676]),.o(intermediate_reg_1[2838])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5675]),.i2(intermediate_reg_0[5674]),.o(intermediate_reg_1[2837]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5673]),.i2(intermediate_reg_0[5672]),.o(intermediate_reg_1[2836]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5671]),.i2(intermediate_reg_0[5670]),.o(intermediate_reg_1[2835])); 
xor_module xor_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5669]),.i2(intermediate_reg_0[5668]),.o(intermediate_reg_1[2834])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5667]),.i2(intermediate_reg_0[5666]),.o(intermediate_reg_1[2833]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5665]),.i2(intermediate_reg_0[5664]),.o(intermediate_reg_1[2832]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5663]),.i2(intermediate_reg_0[5662]),.o(intermediate_reg_1[2831]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5661]),.i2(intermediate_reg_0[5660]),.o(intermediate_reg_1[2830]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5659]),.i2(intermediate_reg_0[5658]),.o(intermediate_reg_1[2829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5657]),.i2(intermediate_reg_0[5656]),.o(intermediate_reg_1[2828]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5655]),.i2(intermediate_reg_0[5654]),.o(intermediate_reg_1[2827])); 
xor_module xor_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5653]),.i2(intermediate_reg_0[5652]),.o(intermediate_reg_1[2826])); 
mux_module mux_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5651]),.i2(intermediate_reg_0[5650]),.o(intermediate_reg_1[2825]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5649]),.i2(intermediate_reg_0[5648]),.o(intermediate_reg_1[2824])); 
xor_module xor_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5647]),.i2(intermediate_reg_0[5646]),.o(intermediate_reg_1[2823])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5645]),.i2(intermediate_reg_0[5644]),.o(intermediate_reg_1[2822]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5643]),.i2(intermediate_reg_0[5642]),.o(intermediate_reg_1[2821])); 
xor_module xor_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5641]),.i2(intermediate_reg_0[5640]),.o(intermediate_reg_1[2820])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5639]),.i2(intermediate_reg_0[5638]),.o(intermediate_reg_1[2819]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5637]),.i2(intermediate_reg_0[5636]),.o(intermediate_reg_1[2818])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5635]),.i2(intermediate_reg_0[5634]),.o(intermediate_reg_1[2817]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5633]),.i2(intermediate_reg_0[5632]),.o(intermediate_reg_1[2816])); 
mux_module mux_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5631]),.i2(intermediate_reg_0[5630]),.o(intermediate_reg_1[2815]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5629]),.i2(intermediate_reg_0[5628]),.o(intermediate_reg_1[2814])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5627]),.i2(intermediate_reg_0[5626]),.o(intermediate_reg_1[2813])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5625]),.i2(intermediate_reg_0[5624]),.o(intermediate_reg_1[2812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5623]),.i2(intermediate_reg_0[5622]),.o(intermediate_reg_1[2811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5621]),.i2(intermediate_reg_0[5620]),.o(intermediate_reg_1[2810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5619]),.i2(intermediate_reg_0[5618]),.o(intermediate_reg_1[2809]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5617]),.i2(intermediate_reg_0[5616]),.o(intermediate_reg_1[2808])); 
xor_module xor_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5615]),.i2(intermediate_reg_0[5614]),.o(intermediate_reg_1[2807])); 
xor_module xor_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5613]),.i2(intermediate_reg_0[5612]),.o(intermediate_reg_1[2806])); 
xor_module xor_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5611]),.i2(intermediate_reg_0[5610]),.o(intermediate_reg_1[2805])); 
xor_module xor_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5609]),.i2(intermediate_reg_0[5608]),.o(intermediate_reg_1[2804])); 
xor_module xor_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5607]),.i2(intermediate_reg_0[5606]),.o(intermediate_reg_1[2803])); 
mux_module mux_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5605]),.i2(intermediate_reg_0[5604]),.o(intermediate_reg_1[2802]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5603]),.i2(intermediate_reg_0[5602]),.o(intermediate_reg_1[2801])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5601]),.i2(intermediate_reg_0[5600]),.o(intermediate_reg_1[2800]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5599]),.i2(intermediate_reg_0[5598]),.o(intermediate_reg_1[2799]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5597]),.i2(intermediate_reg_0[5596]),.o(intermediate_reg_1[2798]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5595]),.i2(intermediate_reg_0[5594]),.o(intermediate_reg_1[2797])); 
mux_module mux_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5593]),.i2(intermediate_reg_0[5592]),.o(intermediate_reg_1[2796]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5591]),.i2(intermediate_reg_0[5590]),.o(intermediate_reg_1[2795])); 
mux_module mux_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5589]),.i2(intermediate_reg_0[5588]),.o(intermediate_reg_1[2794]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5587]),.i2(intermediate_reg_0[5586]),.o(intermediate_reg_1[2793]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5585]),.i2(intermediate_reg_0[5584]),.o(intermediate_reg_1[2792])); 
xor_module xor_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5583]),.i2(intermediate_reg_0[5582]),.o(intermediate_reg_1[2791])); 
xor_module xor_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5581]),.i2(intermediate_reg_0[5580]),.o(intermediate_reg_1[2790])); 
xor_module xor_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5579]),.i2(intermediate_reg_0[5578]),.o(intermediate_reg_1[2789])); 
mux_module mux_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5577]),.i2(intermediate_reg_0[5576]),.o(intermediate_reg_1[2788]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5575]),.i2(intermediate_reg_0[5574]),.o(intermediate_reg_1[2787])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5573]),.i2(intermediate_reg_0[5572]),.o(intermediate_reg_1[2786]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5571]),.i2(intermediate_reg_0[5570]),.o(intermediate_reg_1[2785])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5569]),.i2(intermediate_reg_0[5568]),.o(intermediate_reg_1[2784])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5567]),.i2(intermediate_reg_0[5566]),.o(intermediate_reg_1[2783]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5565]),.i2(intermediate_reg_0[5564]),.o(intermediate_reg_1[2782])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5563]),.i2(intermediate_reg_0[5562]),.o(intermediate_reg_1[2781])); 
mux_module mux_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5561]),.i2(intermediate_reg_0[5560]),.o(intermediate_reg_1[2780]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5559]),.i2(intermediate_reg_0[5558]),.o(intermediate_reg_1[2779])); 
xor_module xor_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5557]),.i2(intermediate_reg_0[5556]),.o(intermediate_reg_1[2778])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5555]),.i2(intermediate_reg_0[5554]),.o(intermediate_reg_1[2777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5553]),.i2(intermediate_reg_0[5552]),.o(intermediate_reg_1[2776]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5551]),.i2(intermediate_reg_0[5550]),.o(intermediate_reg_1[2775])); 
xor_module xor_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5549]),.i2(intermediate_reg_0[5548]),.o(intermediate_reg_1[2774])); 
xor_module xor_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5547]),.i2(intermediate_reg_0[5546]),.o(intermediate_reg_1[2773])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5545]),.i2(intermediate_reg_0[5544]),.o(intermediate_reg_1[2772]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5543]),.i2(intermediate_reg_0[5542]),.o(intermediate_reg_1[2771])); 
xor_module xor_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5541]),.i2(intermediate_reg_0[5540]),.o(intermediate_reg_1[2770])); 
mux_module mux_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5539]),.i2(intermediate_reg_0[5538]),.o(intermediate_reg_1[2769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5537]),.i2(intermediate_reg_0[5536]),.o(intermediate_reg_1[2768]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5535]),.i2(intermediate_reg_0[5534]),.o(intermediate_reg_1[2767])); 
xor_module xor_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5533]),.i2(intermediate_reg_0[5532]),.o(intermediate_reg_1[2766])); 
xor_module xor_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5531]),.i2(intermediate_reg_0[5530]),.o(intermediate_reg_1[2765])); 
xor_module xor_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5529]),.i2(intermediate_reg_0[5528]),.o(intermediate_reg_1[2764])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5527]),.i2(intermediate_reg_0[5526]),.o(intermediate_reg_1[2763])); 
mux_module mux_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5525]),.i2(intermediate_reg_0[5524]),.o(intermediate_reg_1[2762]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5523]),.i2(intermediate_reg_0[5522]),.o(intermediate_reg_1[2761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5521]),.i2(intermediate_reg_0[5520]),.o(intermediate_reg_1[2760]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5519]),.i2(intermediate_reg_0[5518]),.o(intermediate_reg_1[2759]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5517]),.i2(intermediate_reg_0[5516]),.o(intermediate_reg_1[2758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5515]),.i2(intermediate_reg_0[5514]),.o(intermediate_reg_1[2757]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5513]),.i2(intermediate_reg_0[5512]),.o(intermediate_reg_1[2756]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5511]),.i2(intermediate_reg_0[5510]),.o(intermediate_reg_1[2755]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5509]),.i2(intermediate_reg_0[5508]),.o(intermediate_reg_1[2754]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5507]),.i2(intermediate_reg_0[5506]),.o(intermediate_reg_1[2753])); 
xor_module xor_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5505]),.i2(intermediate_reg_0[5504]),.o(intermediate_reg_1[2752])); 
mux_module mux_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5503]),.i2(intermediate_reg_0[5502]),.o(intermediate_reg_1[2751]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5501]),.i2(intermediate_reg_0[5500]),.o(intermediate_reg_1[2750])); 
xor_module xor_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5499]),.i2(intermediate_reg_0[5498]),.o(intermediate_reg_1[2749])); 
xor_module xor_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5497]),.i2(intermediate_reg_0[5496]),.o(intermediate_reg_1[2748])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5495]),.i2(intermediate_reg_0[5494]),.o(intermediate_reg_1[2747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5493]),.i2(intermediate_reg_0[5492]),.o(intermediate_reg_1[2746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5491]),.i2(intermediate_reg_0[5490]),.o(intermediate_reg_1[2745]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5489]),.i2(intermediate_reg_0[5488]),.o(intermediate_reg_1[2744])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5487]),.i2(intermediate_reg_0[5486]),.o(intermediate_reg_1[2743]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5485]),.i2(intermediate_reg_0[5484]),.o(intermediate_reg_1[2742]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5483]),.i2(intermediate_reg_0[5482]),.o(intermediate_reg_1[2741]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5481]),.i2(intermediate_reg_0[5480]),.o(intermediate_reg_1[2740]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5479]),.i2(intermediate_reg_0[5478]),.o(intermediate_reg_1[2739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5477]),.i2(intermediate_reg_0[5476]),.o(intermediate_reg_1[2738]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5475]),.i2(intermediate_reg_0[5474]),.o(intermediate_reg_1[2737]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5473]),.i2(intermediate_reg_0[5472]),.o(intermediate_reg_1[2736]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5471]),.i2(intermediate_reg_0[5470]),.o(intermediate_reg_1[2735]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5469]),.i2(intermediate_reg_0[5468]),.o(intermediate_reg_1[2734]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5467]),.i2(intermediate_reg_0[5466]),.o(intermediate_reg_1[2733]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5465]),.i2(intermediate_reg_0[5464]),.o(intermediate_reg_1[2732])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5463]),.i2(intermediate_reg_0[5462]),.o(intermediate_reg_1[2731]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5461]),.i2(intermediate_reg_0[5460]),.o(intermediate_reg_1[2730])); 
mux_module mux_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5459]),.i2(intermediate_reg_0[5458]),.o(intermediate_reg_1[2729]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5457]),.i2(intermediate_reg_0[5456]),.o(intermediate_reg_1[2728])); 
xor_module xor_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5455]),.i2(intermediate_reg_0[5454]),.o(intermediate_reg_1[2727])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5453]),.i2(intermediate_reg_0[5452]),.o(intermediate_reg_1[2726]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5451]),.i2(intermediate_reg_0[5450]),.o(intermediate_reg_1[2725]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5449]),.i2(intermediate_reg_0[5448]),.o(intermediate_reg_1[2724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5447]),.i2(intermediate_reg_0[5446]),.o(intermediate_reg_1[2723]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5445]),.i2(intermediate_reg_0[5444]),.o(intermediate_reg_1[2722]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5443]),.i2(intermediate_reg_0[5442]),.o(intermediate_reg_1[2721])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5441]),.i2(intermediate_reg_0[5440]),.o(intermediate_reg_1[2720]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5439]),.i2(intermediate_reg_0[5438]),.o(intermediate_reg_1[2719])); 
xor_module xor_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5437]),.i2(intermediate_reg_0[5436]),.o(intermediate_reg_1[2718])); 
xor_module xor_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5435]),.i2(intermediate_reg_0[5434]),.o(intermediate_reg_1[2717])); 
mux_module mux_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5433]),.i2(intermediate_reg_0[5432]),.o(intermediate_reg_1[2716]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5431]),.i2(intermediate_reg_0[5430]),.o(intermediate_reg_1[2715])); 
mux_module mux_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5429]),.i2(intermediate_reg_0[5428]),.o(intermediate_reg_1[2714]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5427]),.i2(intermediate_reg_0[5426]),.o(intermediate_reg_1[2713]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5425]),.i2(intermediate_reg_0[5424]),.o(intermediate_reg_1[2712]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5423]),.i2(intermediate_reg_0[5422]),.o(intermediate_reg_1[2711]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5421]),.i2(intermediate_reg_0[5420]),.o(intermediate_reg_1[2710])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5419]),.i2(intermediate_reg_0[5418]),.o(intermediate_reg_1[2709]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5417]),.i2(intermediate_reg_0[5416]),.o(intermediate_reg_1[2708])); 
xor_module xor_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5415]),.i2(intermediate_reg_0[5414]),.o(intermediate_reg_1[2707])); 
mux_module mux_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5413]),.i2(intermediate_reg_0[5412]),.o(intermediate_reg_1[2706]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5411]),.i2(intermediate_reg_0[5410]),.o(intermediate_reg_1[2705])); 
mux_module mux_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5409]),.i2(intermediate_reg_0[5408]),.o(intermediate_reg_1[2704]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5407]),.i2(intermediate_reg_0[5406]),.o(intermediate_reg_1[2703]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5405]),.i2(intermediate_reg_0[5404]),.o(intermediate_reg_1[2702])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5403]),.i2(intermediate_reg_0[5402]),.o(intermediate_reg_1[2701]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5401]),.i2(intermediate_reg_0[5400]),.o(intermediate_reg_1[2700]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5399]),.i2(intermediate_reg_0[5398]),.o(intermediate_reg_1[2699]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5397]),.i2(intermediate_reg_0[5396]),.o(intermediate_reg_1[2698])); 
mux_module mux_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5395]),.i2(intermediate_reg_0[5394]),.o(intermediate_reg_1[2697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5393]),.i2(intermediate_reg_0[5392]),.o(intermediate_reg_1[2696]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5391]),.i2(intermediate_reg_0[5390]),.o(intermediate_reg_1[2695])); 
mux_module mux_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5389]),.i2(intermediate_reg_0[5388]),.o(intermediate_reg_1[2694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5387]),.i2(intermediate_reg_0[5386]),.o(intermediate_reg_1[2693]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5385]),.i2(intermediate_reg_0[5384]),.o(intermediate_reg_1[2692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5383]),.i2(intermediate_reg_0[5382]),.o(intermediate_reg_1[2691]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5381]),.i2(intermediate_reg_0[5380]),.o(intermediate_reg_1[2690])); 
xor_module xor_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5379]),.i2(intermediate_reg_0[5378]),.o(intermediate_reg_1[2689])); 
xor_module xor_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5377]),.i2(intermediate_reg_0[5376]),.o(intermediate_reg_1[2688])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5375]),.i2(intermediate_reg_0[5374]),.o(intermediate_reg_1[2687]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5373]),.i2(intermediate_reg_0[5372]),.o(intermediate_reg_1[2686])); 
xor_module xor_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5371]),.i2(intermediate_reg_0[5370]),.o(intermediate_reg_1[2685])); 
mux_module mux_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5369]),.i2(intermediate_reg_0[5368]),.o(intermediate_reg_1[2684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5367]),.i2(intermediate_reg_0[5366]),.o(intermediate_reg_1[2683]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5365]),.i2(intermediate_reg_0[5364]),.o(intermediate_reg_1[2682])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5363]),.i2(intermediate_reg_0[5362]),.o(intermediate_reg_1[2681]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5361]),.i2(intermediate_reg_0[5360]),.o(intermediate_reg_1[2680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5359]),.i2(intermediate_reg_0[5358]),.o(intermediate_reg_1[2679]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5357]),.i2(intermediate_reg_0[5356]),.o(intermediate_reg_1[2678])); 
mux_module mux_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5355]),.i2(intermediate_reg_0[5354]),.o(intermediate_reg_1[2677]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5353]),.i2(intermediate_reg_0[5352]),.o(intermediate_reg_1[2676]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5351]),.i2(intermediate_reg_0[5350]),.o(intermediate_reg_1[2675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5349]),.i2(intermediate_reg_0[5348]),.o(intermediate_reg_1[2674]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5347]),.i2(intermediate_reg_0[5346]),.o(intermediate_reg_1[2673])); 
mux_module mux_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5345]),.i2(intermediate_reg_0[5344]),.o(intermediate_reg_1[2672]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5343]),.i2(intermediate_reg_0[5342]),.o(intermediate_reg_1[2671])); 
xor_module xor_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5341]),.i2(intermediate_reg_0[5340]),.o(intermediate_reg_1[2670])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5339]),.i2(intermediate_reg_0[5338]),.o(intermediate_reg_1[2669]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5337]),.i2(intermediate_reg_0[5336]),.o(intermediate_reg_1[2668])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5335]),.i2(intermediate_reg_0[5334]),.o(intermediate_reg_1[2667]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5333]),.i2(intermediate_reg_0[5332]),.o(intermediate_reg_1[2666])); 
mux_module mux_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5331]),.i2(intermediate_reg_0[5330]),.o(intermediate_reg_1[2665]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5329]),.i2(intermediate_reg_0[5328]),.o(intermediate_reg_1[2664]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5327]),.i2(intermediate_reg_0[5326]),.o(intermediate_reg_1[2663])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5325]),.i2(intermediate_reg_0[5324]),.o(intermediate_reg_1[2662])); 
mux_module mux_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5323]),.i2(intermediate_reg_0[5322]),.o(intermediate_reg_1[2661]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5321]),.i2(intermediate_reg_0[5320]),.o(intermediate_reg_1[2660])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5319]),.i2(intermediate_reg_0[5318]),.o(intermediate_reg_1[2659]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5317]),.i2(intermediate_reg_0[5316]),.o(intermediate_reg_1[2658])); 
mux_module mux_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5315]),.i2(intermediate_reg_0[5314]),.o(intermediate_reg_1[2657]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5313]),.i2(intermediate_reg_0[5312]),.o(intermediate_reg_1[2656]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5311]),.i2(intermediate_reg_0[5310]),.o(intermediate_reg_1[2655])); 
xor_module xor_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5309]),.i2(intermediate_reg_0[5308]),.o(intermediate_reg_1[2654])); 
xor_module xor_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5307]),.i2(intermediate_reg_0[5306]),.o(intermediate_reg_1[2653])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5305]),.i2(intermediate_reg_0[5304]),.o(intermediate_reg_1[2652]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5303]),.i2(intermediate_reg_0[5302]),.o(intermediate_reg_1[2651]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5301]),.i2(intermediate_reg_0[5300]),.o(intermediate_reg_1[2650])); 
xor_module xor_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5299]),.i2(intermediate_reg_0[5298]),.o(intermediate_reg_1[2649])); 
xor_module xor_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5297]),.i2(intermediate_reg_0[5296]),.o(intermediate_reg_1[2648])); 
xor_module xor_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5295]),.i2(intermediate_reg_0[5294]),.o(intermediate_reg_1[2647])); 
mux_module mux_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5293]),.i2(intermediate_reg_0[5292]),.o(intermediate_reg_1[2646]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5291]),.i2(intermediate_reg_0[5290]),.o(intermediate_reg_1[2645])); 
xor_module xor_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5289]),.i2(intermediate_reg_0[5288]),.o(intermediate_reg_1[2644])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5287]),.i2(intermediate_reg_0[5286]),.o(intermediate_reg_1[2643]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5285]),.i2(intermediate_reg_0[5284]),.o(intermediate_reg_1[2642])); 
xor_module xor_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5283]),.i2(intermediate_reg_0[5282]),.o(intermediate_reg_1[2641])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5281]),.i2(intermediate_reg_0[5280]),.o(intermediate_reg_1[2640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5279]),.i2(intermediate_reg_0[5278]),.o(intermediate_reg_1[2639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5277]),.i2(intermediate_reg_0[5276]),.o(intermediate_reg_1[2638]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5275]),.i2(intermediate_reg_0[5274]),.o(intermediate_reg_1[2637])); 
xor_module xor_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5273]),.i2(intermediate_reg_0[5272]),.o(intermediate_reg_1[2636])); 
mux_module mux_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5271]),.i2(intermediate_reg_0[5270]),.o(intermediate_reg_1[2635]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5269]),.i2(intermediate_reg_0[5268]),.o(intermediate_reg_1[2634])); 
xor_module xor_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5267]),.i2(intermediate_reg_0[5266]),.o(intermediate_reg_1[2633])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5265]),.i2(intermediate_reg_0[5264]),.o(intermediate_reg_1[2632])); 
xor_module xor_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5263]),.i2(intermediate_reg_0[5262]),.o(intermediate_reg_1[2631])); 
xor_module xor_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5261]),.i2(intermediate_reg_0[5260]),.o(intermediate_reg_1[2630])); 
xor_module xor_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5259]),.i2(intermediate_reg_0[5258]),.o(intermediate_reg_1[2629])); 
xor_module xor_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5257]),.i2(intermediate_reg_0[5256]),.o(intermediate_reg_1[2628])); 
xor_module xor_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5255]),.i2(intermediate_reg_0[5254]),.o(intermediate_reg_1[2627])); 
mux_module mux_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5253]),.i2(intermediate_reg_0[5252]),.o(intermediate_reg_1[2626]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5251]),.i2(intermediate_reg_0[5250]),.o(intermediate_reg_1[2625]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5249]),.i2(intermediate_reg_0[5248]),.o(intermediate_reg_1[2624])); 
mux_module mux_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5247]),.i2(intermediate_reg_0[5246]),.o(intermediate_reg_1[2623]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5245]),.i2(intermediate_reg_0[5244]),.o(intermediate_reg_1[2622]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5243]),.i2(intermediate_reg_0[5242]),.o(intermediate_reg_1[2621]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5241]),.i2(intermediate_reg_0[5240]),.o(intermediate_reg_1[2620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5239]),.i2(intermediate_reg_0[5238]),.o(intermediate_reg_1[2619]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5237]),.i2(intermediate_reg_0[5236]),.o(intermediate_reg_1[2618])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5235]),.i2(intermediate_reg_0[5234]),.o(intermediate_reg_1[2617]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5233]),.i2(intermediate_reg_0[5232]),.o(intermediate_reg_1[2616])); 
mux_module mux_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5231]),.i2(intermediate_reg_0[5230]),.o(intermediate_reg_1[2615]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5229]),.i2(intermediate_reg_0[5228]),.o(intermediate_reg_1[2614])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5227]),.i2(intermediate_reg_0[5226]),.o(intermediate_reg_1[2613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5225]),.i2(intermediate_reg_0[5224]),.o(intermediate_reg_1[2612]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5223]),.i2(intermediate_reg_0[5222]),.o(intermediate_reg_1[2611]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5221]),.i2(intermediate_reg_0[5220]),.o(intermediate_reg_1[2610])); 
xor_module xor_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5219]),.i2(intermediate_reg_0[5218]),.o(intermediate_reg_1[2609])); 
mux_module mux_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5217]),.i2(intermediate_reg_0[5216]),.o(intermediate_reg_1[2608]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5215]),.i2(intermediate_reg_0[5214]),.o(intermediate_reg_1[2607])); 
xor_module xor_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5213]),.i2(intermediate_reg_0[5212]),.o(intermediate_reg_1[2606])); 
xor_module xor_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5211]),.i2(intermediate_reg_0[5210]),.o(intermediate_reg_1[2605])); 
xor_module xor_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5209]),.i2(intermediate_reg_0[5208]),.o(intermediate_reg_1[2604])); 
mux_module mux_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5207]),.i2(intermediate_reg_0[5206]),.o(intermediate_reg_1[2603]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5205]),.i2(intermediate_reg_0[5204]),.o(intermediate_reg_1[2602])); 
mux_module mux_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5203]),.i2(intermediate_reg_0[5202]),.o(intermediate_reg_1[2601]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5201]),.i2(intermediate_reg_0[5200]),.o(intermediate_reg_1[2600])); 
xor_module xor_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5199]),.i2(intermediate_reg_0[5198]),.o(intermediate_reg_1[2599])); 
xor_module xor_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5197]),.i2(intermediate_reg_0[5196]),.o(intermediate_reg_1[2598])); 
xor_module xor_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5195]),.i2(intermediate_reg_0[5194]),.o(intermediate_reg_1[2597])); 
xor_module xor_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5193]),.i2(intermediate_reg_0[5192]),.o(intermediate_reg_1[2596])); 
xor_module xor_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5191]),.i2(intermediate_reg_0[5190]),.o(intermediate_reg_1[2595])); 
mux_module mux_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5189]),.i2(intermediate_reg_0[5188]),.o(intermediate_reg_1[2594]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5187]),.i2(intermediate_reg_0[5186]),.o(intermediate_reg_1[2593]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5185]),.i2(intermediate_reg_0[5184]),.o(intermediate_reg_1[2592])); 
mux_module mux_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5183]),.i2(intermediate_reg_0[5182]),.o(intermediate_reg_1[2591]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5181]),.i2(intermediate_reg_0[5180]),.o(intermediate_reg_1[2590])); 
mux_module mux_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5179]),.i2(intermediate_reg_0[5178]),.o(intermediate_reg_1[2589]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5177]),.i2(intermediate_reg_0[5176]),.o(intermediate_reg_1[2588])); 
mux_module mux_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5175]),.i2(intermediate_reg_0[5174]),.o(intermediate_reg_1[2587]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5173]),.i2(intermediate_reg_0[5172]),.o(intermediate_reg_1[2586])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5171]),.i2(intermediate_reg_0[5170]),.o(intermediate_reg_1[2585]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5169]),.i2(intermediate_reg_0[5168]),.o(intermediate_reg_1[2584])); 
xor_module xor_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5167]),.i2(intermediate_reg_0[5166]),.o(intermediate_reg_1[2583])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5165]),.i2(intermediate_reg_0[5164]),.o(intermediate_reg_1[2582])); 
mux_module mux_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5163]),.i2(intermediate_reg_0[5162]),.o(intermediate_reg_1[2581]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5161]),.i2(intermediate_reg_0[5160]),.o(intermediate_reg_1[2580]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5159]),.i2(intermediate_reg_0[5158]),.o(intermediate_reg_1[2579]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5157]),.i2(intermediate_reg_0[5156]),.o(intermediate_reg_1[2578])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5155]),.i2(intermediate_reg_0[5154]),.o(intermediate_reg_1[2577]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5153]),.i2(intermediate_reg_0[5152]),.o(intermediate_reg_1[2576]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5151]),.i2(intermediate_reg_0[5150]),.o(intermediate_reg_1[2575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5149]),.i2(intermediate_reg_0[5148]),.o(intermediate_reg_1[2574]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5147]),.i2(intermediate_reg_0[5146]),.o(intermediate_reg_1[2573])); 
xor_module xor_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5145]),.i2(intermediate_reg_0[5144]),.o(intermediate_reg_1[2572])); 
xor_module xor_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5143]),.i2(intermediate_reg_0[5142]),.o(intermediate_reg_1[2571])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5141]),.i2(intermediate_reg_0[5140]),.o(intermediate_reg_1[2570]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5139]),.i2(intermediate_reg_0[5138]),.o(intermediate_reg_1[2569])); 
xor_module xor_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5137]),.i2(intermediate_reg_0[5136]),.o(intermediate_reg_1[2568])); 
xor_module xor_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5135]),.i2(intermediate_reg_0[5134]),.o(intermediate_reg_1[2567])); 
xor_module xor_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5133]),.i2(intermediate_reg_0[5132]),.o(intermediate_reg_1[2566])); 
xor_module xor_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5131]),.i2(intermediate_reg_0[5130]),.o(intermediate_reg_1[2565])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5129]),.i2(intermediate_reg_0[5128]),.o(intermediate_reg_1[2564]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5127]),.i2(intermediate_reg_0[5126]),.o(intermediate_reg_1[2563]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5125]),.i2(intermediate_reg_0[5124]),.o(intermediate_reg_1[2562])); 
xor_module xor_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5123]),.i2(intermediate_reg_0[5122]),.o(intermediate_reg_1[2561])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5121]),.i2(intermediate_reg_0[5120]),.o(intermediate_reg_1[2560]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5119]),.i2(intermediate_reg_0[5118]),.o(intermediate_reg_1[2559])); 
xor_module xor_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5117]),.i2(intermediate_reg_0[5116]),.o(intermediate_reg_1[2558])); 
mux_module mux_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5115]),.i2(intermediate_reg_0[5114]),.o(intermediate_reg_1[2557]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5113]),.i2(intermediate_reg_0[5112]),.o(intermediate_reg_1[2556])); 
mux_module mux_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5111]),.i2(intermediate_reg_0[5110]),.o(intermediate_reg_1[2555]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5109]),.i2(intermediate_reg_0[5108]),.o(intermediate_reg_1[2554])); 
mux_module mux_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5107]),.i2(intermediate_reg_0[5106]),.o(intermediate_reg_1[2553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5105]),.i2(intermediate_reg_0[5104]),.o(intermediate_reg_1[2552]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5103]),.i2(intermediate_reg_0[5102]),.o(intermediate_reg_1[2551]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5101]),.i2(intermediate_reg_0[5100]),.o(intermediate_reg_1[2550]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5099]),.i2(intermediate_reg_0[5098]),.o(intermediate_reg_1[2549]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5097]),.i2(intermediate_reg_0[5096]),.o(intermediate_reg_1[2548])); 
mux_module mux_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5095]),.i2(intermediate_reg_0[5094]),.o(intermediate_reg_1[2547]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5093]),.i2(intermediate_reg_0[5092]),.o(intermediate_reg_1[2546]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5091]),.i2(intermediate_reg_0[5090]),.o(intermediate_reg_1[2545])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5089]),.i2(intermediate_reg_0[5088]),.o(intermediate_reg_1[2544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5087]),.i2(intermediate_reg_0[5086]),.o(intermediate_reg_1[2543]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5085]),.i2(intermediate_reg_0[5084]),.o(intermediate_reg_1[2542])); 
xor_module xor_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5083]),.i2(intermediate_reg_0[5082]),.o(intermediate_reg_1[2541])); 
xor_module xor_module_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5081]),.i2(intermediate_reg_0[5080]),.o(intermediate_reg_1[2540])); 
xor_module xor_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5079]),.i2(intermediate_reg_0[5078]),.o(intermediate_reg_1[2539])); 
xor_module xor_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5077]),.i2(intermediate_reg_0[5076]),.o(intermediate_reg_1[2538])); 
mux_module mux_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5075]),.i2(intermediate_reg_0[5074]),.o(intermediate_reg_1[2537]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5073]),.i2(intermediate_reg_0[5072]),.o(intermediate_reg_1[2536])); 
xor_module xor_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5071]),.i2(intermediate_reg_0[5070]),.o(intermediate_reg_1[2535])); 
xor_module xor_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5069]),.i2(intermediate_reg_0[5068]),.o(intermediate_reg_1[2534])); 
xor_module xor_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5067]),.i2(intermediate_reg_0[5066]),.o(intermediate_reg_1[2533])); 
xor_module xor_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5065]),.i2(intermediate_reg_0[5064]),.o(intermediate_reg_1[2532])); 
xor_module xor_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5063]),.i2(intermediate_reg_0[5062]),.o(intermediate_reg_1[2531])); 
xor_module xor_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5061]),.i2(intermediate_reg_0[5060]),.o(intermediate_reg_1[2530])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5059]),.i2(intermediate_reg_0[5058]),.o(intermediate_reg_1[2529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5057]),.i2(intermediate_reg_0[5056]),.o(intermediate_reg_1[2528]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5055]),.i2(intermediate_reg_0[5054]),.o(intermediate_reg_1[2527])); 
xor_module xor_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5053]),.i2(intermediate_reg_0[5052]),.o(intermediate_reg_1[2526])); 
mux_module mux_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5051]),.i2(intermediate_reg_0[5050]),.o(intermediate_reg_1[2525]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5049]),.i2(intermediate_reg_0[5048]),.o(intermediate_reg_1[2524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5047]),.i2(intermediate_reg_0[5046]),.o(intermediate_reg_1[2523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5045]),.i2(intermediate_reg_0[5044]),.o(intermediate_reg_1[2522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5043]),.i2(intermediate_reg_0[5042]),.o(intermediate_reg_1[2521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5041]),.i2(intermediate_reg_0[5040]),.o(intermediate_reg_1[2520]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5039]),.i2(intermediate_reg_0[5038]),.o(intermediate_reg_1[2519])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5037]),.i2(intermediate_reg_0[5036]),.o(intermediate_reg_1[2518])); 
xor_module xor_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5035]),.i2(intermediate_reg_0[5034]),.o(intermediate_reg_1[2517])); 
mux_module mux_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5033]),.i2(intermediate_reg_0[5032]),.o(intermediate_reg_1[2516]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5031]),.i2(intermediate_reg_0[5030]),.o(intermediate_reg_1[2515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5029]),.i2(intermediate_reg_0[5028]),.o(intermediate_reg_1[2514]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5027]),.i2(intermediate_reg_0[5026]),.o(intermediate_reg_1[2513]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5025]),.i2(intermediate_reg_0[5024]),.o(intermediate_reg_1[2512])); 
xor_module xor_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5023]),.i2(intermediate_reg_0[5022]),.o(intermediate_reg_1[2511])); 
xor_module xor_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5021]),.i2(intermediate_reg_0[5020]),.o(intermediate_reg_1[2510])); 
xor_module xor_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5019]),.i2(intermediate_reg_0[5018]),.o(intermediate_reg_1[2509])); 
xor_module xor_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5017]),.i2(intermediate_reg_0[5016]),.o(intermediate_reg_1[2508])); 
mux_module mux_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5015]),.i2(intermediate_reg_0[5014]),.o(intermediate_reg_1[2507]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5013]),.i2(intermediate_reg_0[5012]),.o(intermediate_reg_1[2506]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5011]),.i2(intermediate_reg_0[5010]),.o(intermediate_reg_1[2505]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5009]),.i2(intermediate_reg_0[5008]),.o(intermediate_reg_1[2504])); 
mux_module mux_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5007]),.i2(intermediate_reg_0[5006]),.o(intermediate_reg_1[2503]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5005]),.i2(intermediate_reg_0[5004]),.o(intermediate_reg_1[2502]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5003]),.i2(intermediate_reg_0[5002]),.o(intermediate_reg_1[2501]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5001]),.i2(intermediate_reg_0[5000]),.o(intermediate_reg_1[2500])); 
xor_module xor_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4999]),.i2(intermediate_reg_0[4998]),.o(intermediate_reg_1[2499])); 
xor_module xor_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4997]),.i2(intermediate_reg_0[4996]),.o(intermediate_reg_1[2498])); 
xor_module xor_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4995]),.i2(intermediate_reg_0[4994]),.o(intermediate_reg_1[2497])); 
xor_module xor_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4993]),.i2(intermediate_reg_0[4992]),.o(intermediate_reg_1[2496])); 
xor_module xor_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4991]),.i2(intermediate_reg_0[4990]),.o(intermediate_reg_1[2495])); 
mux_module mux_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4989]),.i2(intermediate_reg_0[4988]),.o(intermediate_reg_1[2494]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4987]),.i2(intermediate_reg_0[4986]),.o(intermediate_reg_1[2493]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4985]),.i2(intermediate_reg_0[4984]),.o(intermediate_reg_1[2492])); 
xor_module xor_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4983]),.i2(intermediate_reg_0[4982]),.o(intermediate_reg_1[2491])); 
xor_module xor_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4981]),.i2(intermediate_reg_0[4980]),.o(intermediate_reg_1[2490])); 
mux_module mux_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4979]),.i2(intermediate_reg_0[4978]),.o(intermediate_reg_1[2489]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4977]),.i2(intermediate_reg_0[4976]),.o(intermediate_reg_1[2488])); 
xor_module xor_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4975]),.i2(intermediate_reg_0[4974]),.o(intermediate_reg_1[2487])); 
xor_module xor_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4973]),.i2(intermediate_reg_0[4972]),.o(intermediate_reg_1[2486])); 
xor_module xor_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4971]),.i2(intermediate_reg_0[4970]),.o(intermediate_reg_1[2485])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4969]),.i2(intermediate_reg_0[4968]),.o(intermediate_reg_1[2484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4967]),.i2(intermediate_reg_0[4966]),.o(intermediate_reg_1[2483]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4965]),.i2(intermediate_reg_0[4964]),.o(intermediate_reg_1[2482]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4963]),.i2(intermediate_reg_0[4962]),.o(intermediate_reg_1[2481])); 
mux_module mux_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4961]),.i2(intermediate_reg_0[4960]),.o(intermediate_reg_1[2480]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4959]),.i2(intermediate_reg_0[4958]),.o(intermediate_reg_1[2479]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4957]),.i2(intermediate_reg_0[4956]),.o(intermediate_reg_1[2478])); 
mux_module mux_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4955]),.i2(intermediate_reg_0[4954]),.o(intermediate_reg_1[2477]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4953]),.i2(intermediate_reg_0[4952]),.o(intermediate_reg_1[2476])); 
xor_module xor_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4951]),.i2(intermediate_reg_0[4950]),.o(intermediate_reg_1[2475])); 
xor_module xor_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4949]),.i2(intermediate_reg_0[4948]),.o(intermediate_reg_1[2474])); 
xor_module xor_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4947]),.i2(intermediate_reg_0[4946]),.o(intermediate_reg_1[2473])); 
xor_module xor_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4945]),.i2(intermediate_reg_0[4944]),.o(intermediate_reg_1[2472])); 
mux_module mux_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4943]),.i2(intermediate_reg_0[4942]),.o(intermediate_reg_1[2471]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4941]),.i2(intermediate_reg_0[4940]),.o(intermediate_reg_1[2470]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4939]),.i2(intermediate_reg_0[4938]),.o(intermediate_reg_1[2469])); 
mux_module mux_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4937]),.i2(intermediate_reg_0[4936]),.o(intermediate_reg_1[2468]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4935]),.i2(intermediate_reg_0[4934]),.o(intermediate_reg_1[2467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4933]),.i2(intermediate_reg_0[4932]),.o(intermediate_reg_1[2466]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4931]),.i2(intermediate_reg_0[4930]),.o(intermediate_reg_1[2465])); 
mux_module mux_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4929]),.i2(intermediate_reg_0[4928]),.o(intermediate_reg_1[2464]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4927]),.i2(intermediate_reg_0[4926]),.o(intermediate_reg_1[2463])); 
mux_module mux_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4925]),.i2(intermediate_reg_0[4924]),.o(intermediate_reg_1[2462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4923]),.i2(intermediate_reg_0[4922]),.o(intermediate_reg_1[2461]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4921]),.i2(intermediate_reg_0[4920]),.o(intermediate_reg_1[2460]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4919]),.i2(intermediate_reg_0[4918]),.o(intermediate_reg_1[2459])); 
mux_module mux_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4917]),.i2(intermediate_reg_0[4916]),.o(intermediate_reg_1[2458]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4915]),.i2(intermediate_reg_0[4914]),.o(intermediate_reg_1[2457])); 
xor_module xor_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4913]),.i2(intermediate_reg_0[4912]),.o(intermediate_reg_1[2456])); 
mux_module mux_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4911]),.i2(intermediate_reg_0[4910]),.o(intermediate_reg_1[2455]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4909]),.i2(intermediate_reg_0[4908]),.o(intermediate_reg_1[2454])); 
xor_module xor_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4907]),.i2(intermediate_reg_0[4906]),.o(intermediate_reg_1[2453])); 
mux_module mux_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4905]),.i2(intermediate_reg_0[4904]),.o(intermediate_reg_1[2452]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4903]),.i2(intermediate_reg_0[4902]),.o(intermediate_reg_1[2451]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4901]),.i2(intermediate_reg_0[4900]),.o(intermediate_reg_1[2450])); 
mux_module mux_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4899]),.i2(intermediate_reg_0[4898]),.o(intermediate_reg_1[2449]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4897]),.i2(intermediate_reg_0[4896]),.o(intermediate_reg_1[2448]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4895]),.i2(intermediate_reg_0[4894]),.o(intermediate_reg_1[2447])); 
mux_module mux_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4893]),.i2(intermediate_reg_0[4892]),.o(intermediate_reg_1[2446]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4891]),.i2(intermediate_reg_0[4890]),.o(intermediate_reg_1[2445])); 
xor_module xor_module_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4889]),.i2(intermediate_reg_0[4888]),.o(intermediate_reg_1[2444])); 
xor_module xor_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4887]),.i2(intermediate_reg_0[4886]),.o(intermediate_reg_1[2443])); 
mux_module mux_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4885]),.i2(intermediate_reg_0[4884]),.o(intermediate_reg_1[2442]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4883]),.i2(intermediate_reg_0[4882]),.o(intermediate_reg_1[2441]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4881]),.i2(intermediate_reg_0[4880]),.o(intermediate_reg_1[2440])); 
mux_module mux_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4879]),.i2(intermediate_reg_0[4878]),.o(intermediate_reg_1[2439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4877]),.i2(intermediate_reg_0[4876]),.o(intermediate_reg_1[2438]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4875]),.i2(intermediate_reg_0[4874]),.o(intermediate_reg_1[2437]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4873]),.i2(intermediate_reg_0[4872]),.o(intermediate_reg_1[2436])); 
xor_module xor_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4871]),.i2(intermediate_reg_0[4870]),.o(intermediate_reg_1[2435])); 
mux_module mux_module_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4869]),.i2(intermediate_reg_0[4868]),.o(intermediate_reg_1[2434]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4867]),.i2(intermediate_reg_0[4866]),.o(intermediate_reg_1[2433])); 
mux_module mux_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4865]),.i2(intermediate_reg_0[4864]),.o(intermediate_reg_1[2432]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4863]),.i2(intermediate_reg_0[4862]),.o(intermediate_reg_1[2431])); 
mux_module mux_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4861]),.i2(intermediate_reg_0[4860]),.o(intermediate_reg_1[2430]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4859]),.i2(intermediate_reg_0[4858]),.o(intermediate_reg_1[2429]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4857]),.i2(intermediate_reg_0[4856]),.o(intermediate_reg_1[2428]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4855]),.i2(intermediate_reg_0[4854]),.o(intermediate_reg_1[2427])); 
mux_module mux_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4853]),.i2(intermediate_reg_0[4852]),.o(intermediate_reg_1[2426]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4851]),.i2(intermediate_reg_0[4850]),.o(intermediate_reg_1[2425])); 
mux_module mux_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4849]),.i2(intermediate_reg_0[4848]),.o(intermediate_reg_1[2424]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4847]),.i2(intermediate_reg_0[4846]),.o(intermediate_reg_1[2423])); 
xor_module xor_module_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4845]),.i2(intermediate_reg_0[4844]),.o(intermediate_reg_1[2422])); 
xor_module xor_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4843]),.i2(intermediate_reg_0[4842]),.o(intermediate_reg_1[2421])); 
xor_module xor_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4841]),.i2(intermediate_reg_0[4840]),.o(intermediate_reg_1[2420])); 
mux_module mux_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4839]),.i2(intermediate_reg_0[4838]),.o(intermediate_reg_1[2419]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4837]),.i2(intermediate_reg_0[4836]),.o(intermediate_reg_1[2418])); 
mux_module mux_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4835]),.i2(intermediate_reg_0[4834]),.o(intermediate_reg_1[2417]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4833]),.i2(intermediate_reg_0[4832]),.o(intermediate_reg_1[2416])); 
xor_module xor_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4831]),.i2(intermediate_reg_0[4830]),.o(intermediate_reg_1[2415])); 
xor_module xor_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4829]),.i2(intermediate_reg_0[4828]),.o(intermediate_reg_1[2414])); 
mux_module mux_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4827]),.i2(intermediate_reg_0[4826]),.o(intermediate_reg_1[2413]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4825]),.i2(intermediate_reg_0[4824]),.o(intermediate_reg_1[2412])); 
mux_module mux_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4823]),.i2(intermediate_reg_0[4822]),.o(intermediate_reg_1[2411]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4821]),.i2(intermediate_reg_0[4820]),.o(intermediate_reg_1[2410])); 
xor_module xor_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4819]),.i2(intermediate_reg_0[4818]),.o(intermediate_reg_1[2409])); 
mux_module mux_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4817]),.i2(intermediate_reg_0[4816]),.o(intermediate_reg_1[2408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4815]),.i2(intermediate_reg_0[4814]),.o(intermediate_reg_1[2407]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4813]),.i2(intermediate_reg_0[4812]),.o(intermediate_reg_1[2406]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4811]),.i2(intermediate_reg_0[4810]),.o(intermediate_reg_1[2405])); 
xor_module xor_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4809]),.i2(intermediate_reg_0[4808]),.o(intermediate_reg_1[2404])); 
mux_module mux_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4807]),.i2(intermediate_reg_0[4806]),.o(intermediate_reg_1[2403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4805]),.i2(intermediate_reg_0[4804]),.o(intermediate_reg_1[2402]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4803]),.i2(intermediate_reg_0[4802]),.o(intermediate_reg_1[2401])); 
mux_module mux_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4801]),.i2(intermediate_reg_0[4800]),.o(intermediate_reg_1[2400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4799]),.i2(intermediate_reg_0[4798]),.o(intermediate_reg_1[2399]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4797]),.i2(intermediate_reg_0[4796]),.o(intermediate_reg_1[2398]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4795]),.i2(intermediate_reg_0[4794]),.o(intermediate_reg_1[2397])); 
mux_module mux_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4793]),.i2(intermediate_reg_0[4792]),.o(intermediate_reg_1[2396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4791]),.i2(intermediate_reg_0[4790]),.o(intermediate_reg_1[2395])); 
mux_module mux_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4789]),.i2(intermediate_reg_0[4788]),.o(intermediate_reg_1[2394]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4787]),.i2(intermediate_reg_0[4786]),.o(intermediate_reg_1[2393]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4785]),.i2(intermediate_reg_0[4784]),.o(intermediate_reg_1[2392]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4783]),.i2(intermediate_reg_0[4782]),.o(intermediate_reg_1[2391]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4781]),.i2(intermediate_reg_0[4780]),.o(intermediate_reg_1[2390]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4779]),.i2(intermediate_reg_0[4778]),.o(intermediate_reg_1[2389]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4777]),.i2(intermediate_reg_0[4776]),.o(intermediate_reg_1[2388])); 
mux_module mux_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4775]),.i2(intermediate_reg_0[4774]),.o(intermediate_reg_1[2387]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4773]),.i2(intermediate_reg_0[4772]),.o(intermediate_reg_1[2386])); 
xor_module xor_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4771]),.i2(intermediate_reg_0[4770]),.o(intermediate_reg_1[2385])); 
mux_module mux_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4769]),.i2(intermediate_reg_0[4768]),.o(intermediate_reg_1[2384]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4767]),.i2(intermediate_reg_0[4766]),.o(intermediate_reg_1[2383]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4765]),.i2(intermediate_reg_0[4764]),.o(intermediate_reg_1[2382]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4763]),.i2(intermediate_reg_0[4762]),.o(intermediate_reg_1[2381])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4761]),.i2(intermediate_reg_0[4760]),.o(intermediate_reg_1[2380]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4759]),.i2(intermediate_reg_0[4758]),.o(intermediate_reg_1[2379])); 
mux_module mux_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4757]),.i2(intermediate_reg_0[4756]),.o(intermediate_reg_1[2378]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4755]),.i2(intermediate_reg_0[4754]),.o(intermediate_reg_1[2377])); 
mux_module mux_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4753]),.i2(intermediate_reg_0[4752]),.o(intermediate_reg_1[2376]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4751]),.i2(intermediate_reg_0[4750]),.o(intermediate_reg_1[2375]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4749]),.i2(intermediate_reg_0[4748]),.o(intermediate_reg_1[2374])); 
xor_module xor_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4747]),.i2(intermediate_reg_0[4746]),.o(intermediate_reg_1[2373])); 
mux_module mux_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4745]),.i2(intermediate_reg_0[4744]),.o(intermediate_reg_1[2372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4743]),.i2(intermediate_reg_0[4742]),.o(intermediate_reg_1[2371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4741]),.i2(intermediate_reg_0[4740]),.o(intermediate_reg_1[2370]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4739]),.i2(intermediate_reg_0[4738]),.o(intermediate_reg_1[2369]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4737]),.i2(intermediate_reg_0[4736]),.o(intermediate_reg_1[2368])); 
xor_module xor_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4735]),.i2(intermediate_reg_0[4734]),.o(intermediate_reg_1[2367])); 
xor_module xor_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4733]),.i2(intermediate_reg_0[4732]),.o(intermediate_reg_1[2366])); 
xor_module xor_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4731]),.i2(intermediate_reg_0[4730]),.o(intermediate_reg_1[2365])); 
mux_module mux_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4729]),.i2(intermediate_reg_0[4728]),.o(intermediate_reg_1[2364]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4727]),.i2(intermediate_reg_0[4726]),.o(intermediate_reg_1[2363])); 
mux_module mux_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4725]),.i2(intermediate_reg_0[4724]),.o(intermediate_reg_1[2362]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4723]),.i2(intermediate_reg_0[4722]),.o(intermediate_reg_1[2361]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4721]),.i2(intermediate_reg_0[4720]),.o(intermediate_reg_1[2360])); 
xor_module xor_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4719]),.i2(intermediate_reg_0[4718]),.o(intermediate_reg_1[2359])); 
mux_module mux_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4717]),.i2(intermediate_reg_0[4716]),.o(intermediate_reg_1[2358]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4715]),.i2(intermediate_reg_0[4714]),.o(intermediate_reg_1[2357]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4713]),.i2(intermediate_reg_0[4712]),.o(intermediate_reg_1[2356])); 
xor_module xor_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4711]),.i2(intermediate_reg_0[4710]),.o(intermediate_reg_1[2355])); 
mux_module mux_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4709]),.i2(intermediate_reg_0[4708]),.o(intermediate_reg_1[2354]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4707]),.i2(intermediate_reg_0[4706]),.o(intermediate_reg_1[2353])); 
mux_module mux_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4705]),.i2(intermediate_reg_0[4704]),.o(intermediate_reg_1[2352]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4703]),.i2(intermediate_reg_0[4702]),.o(intermediate_reg_1[2351])); 
xor_module xor_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4701]),.i2(intermediate_reg_0[4700]),.o(intermediate_reg_1[2350])); 
mux_module mux_module_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4699]),.i2(intermediate_reg_0[4698]),.o(intermediate_reg_1[2349]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4697]),.i2(intermediate_reg_0[4696]),.o(intermediate_reg_1[2348])); 
xor_module xor_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4695]),.i2(intermediate_reg_0[4694]),.o(intermediate_reg_1[2347])); 
mux_module mux_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4693]),.i2(intermediate_reg_0[4692]),.o(intermediate_reg_1[2346]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4691]),.i2(intermediate_reg_0[4690]),.o(intermediate_reg_1[2345])); 
mux_module mux_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4689]),.i2(intermediate_reg_0[4688]),.o(intermediate_reg_1[2344]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4687]),.i2(intermediate_reg_0[4686]),.o(intermediate_reg_1[2343]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4685]),.i2(intermediate_reg_0[4684]),.o(intermediate_reg_1[2342])); 
xor_module xor_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4683]),.i2(intermediate_reg_0[4682]),.o(intermediate_reg_1[2341])); 
mux_module mux_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4681]),.i2(intermediate_reg_0[4680]),.o(intermediate_reg_1[2340]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4679]),.i2(intermediate_reg_0[4678]),.o(intermediate_reg_1[2339]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4677]),.i2(intermediate_reg_0[4676]),.o(intermediate_reg_1[2338])); 
mux_module mux_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4675]),.i2(intermediate_reg_0[4674]),.o(intermediate_reg_1[2337]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4673]),.i2(intermediate_reg_0[4672]),.o(intermediate_reg_1[2336])); 
mux_module mux_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4671]),.i2(intermediate_reg_0[4670]),.o(intermediate_reg_1[2335]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4669]),.i2(intermediate_reg_0[4668]),.o(intermediate_reg_1[2334])); 
mux_module mux_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4667]),.i2(intermediate_reg_0[4666]),.o(intermediate_reg_1[2333]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4665]),.i2(intermediate_reg_0[4664]),.o(intermediate_reg_1[2332])); 
xor_module xor_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4663]),.i2(intermediate_reg_0[4662]),.o(intermediate_reg_1[2331])); 
xor_module xor_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4661]),.i2(intermediate_reg_0[4660]),.o(intermediate_reg_1[2330])); 
mux_module mux_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4659]),.i2(intermediate_reg_0[4658]),.o(intermediate_reg_1[2329]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4657]),.i2(intermediate_reg_0[4656]),.o(intermediate_reg_1[2328])); 
mux_module mux_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4655]),.i2(intermediate_reg_0[4654]),.o(intermediate_reg_1[2327]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4653]),.i2(intermediate_reg_0[4652]),.o(intermediate_reg_1[2326]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4651]),.i2(intermediate_reg_0[4650]),.o(intermediate_reg_1[2325])); 
mux_module mux_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4649]),.i2(intermediate_reg_0[4648]),.o(intermediate_reg_1[2324]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4647]),.i2(intermediate_reg_0[4646]),.o(intermediate_reg_1[2323])); 
xor_module xor_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4645]),.i2(intermediate_reg_0[4644]),.o(intermediate_reg_1[2322])); 
mux_module mux_module_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4643]),.i2(intermediate_reg_0[4642]),.o(intermediate_reg_1[2321]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4641]),.i2(intermediate_reg_0[4640]),.o(intermediate_reg_1[2320]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4639]),.i2(intermediate_reg_0[4638]),.o(intermediate_reg_1[2319])); 
mux_module mux_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4637]),.i2(intermediate_reg_0[4636]),.o(intermediate_reg_1[2318]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4635]),.i2(intermediate_reg_0[4634]),.o(intermediate_reg_1[2317])); 
xor_module xor_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4633]),.i2(intermediate_reg_0[4632]),.o(intermediate_reg_1[2316])); 
mux_module mux_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4631]),.i2(intermediate_reg_0[4630]),.o(intermediate_reg_1[2315]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4629]),.i2(intermediate_reg_0[4628]),.o(intermediate_reg_1[2314]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4627]),.i2(intermediate_reg_0[4626]),.o(intermediate_reg_1[2313]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4625]),.i2(intermediate_reg_0[4624]),.o(intermediate_reg_1[2312])); 
xor_module xor_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4623]),.i2(intermediate_reg_0[4622]),.o(intermediate_reg_1[2311])); 
xor_module xor_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4621]),.i2(intermediate_reg_0[4620]),.o(intermediate_reg_1[2310])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4619]),.i2(intermediate_reg_0[4618]),.o(intermediate_reg_1[2309]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4617]),.i2(intermediate_reg_0[4616]),.o(intermediate_reg_1[2308])); 
xor_module xor_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4615]),.i2(intermediate_reg_0[4614]),.o(intermediate_reg_1[2307])); 
xor_module xor_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4613]),.i2(intermediate_reg_0[4612]),.o(intermediate_reg_1[2306])); 
mux_module mux_module_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4611]),.i2(intermediate_reg_0[4610]),.o(intermediate_reg_1[2305]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4609]),.i2(intermediate_reg_0[4608]),.o(intermediate_reg_1[2304])); 
mux_module mux_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4607]),.i2(intermediate_reg_0[4606]),.o(intermediate_reg_1[2303]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4605]),.i2(intermediate_reg_0[4604]),.o(intermediate_reg_1[2302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4603]),.i2(intermediate_reg_0[4602]),.o(intermediate_reg_1[2301]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4601]),.i2(intermediate_reg_0[4600]),.o(intermediate_reg_1[2300]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4599]),.i2(intermediate_reg_0[4598]),.o(intermediate_reg_1[2299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4597]),.i2(intermediate_reg_0[4596]),.o(intermediate_reg_1[2298]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4595]),.i2(intermediate_reg_0[4594]),.o(intermediate_reg_1[2297])); 
xor_module xor_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4593]),.i2(intermediate_reg_0[4592]),.o(intermediate_reg_1[2296])); 
xor_module xor_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4591]),.i2(intermediate_reg_0[4590]),.o(intermediate_reg_1[2295])); 
xor_module xor_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4589]),.i2(intermediate_reg_0[4588]),.o(intermediate_reg_1[2294])); 
xor_module xor_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4587]),.i2(intermediate_reg_0[4586]),.o(intermediate_reg_1[2293])); 
xor_module xor_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4585]),.i2(intermediate_reg_0[4584]),.o(intermediate_reg_1[2292])); 
xor_module xor_module_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4583]),.i2(intermediate_reg_0[4582]),.o(intermediate_reg_1[2291])); 
mux_module mux_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4581]),.i2(intermediate_reg_0[4580]),.o(intermediate_reg_1[2290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4579]),.i2(intermediate_reg_0[4578]),.o(intermediate_reg_1[2289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4577]),.i2(intermediate_reg_0[4576]),.o(intermediate_reg_1[2288]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4575]),.i2(intermediate_reg_0[4574]),.o(intermediate_reg_1[2287]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4573]),.i2(intermediate_reg_0[4572]),.o(intermediate_reg_1[2286])); 
mux_module mux_module_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4571]),.i2(intermediate_reg_0[4570]),.o(intermediate_reg_1[2285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4569]),.i2(intermediate_reg_0[4568]),.o(intermediate_reg_1[2284]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4567]),.i2(intermediate_reg_0[4566]),.o(intermediate_reg_1[2283])); 
mux_module mux_module_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4565]),.i2(intermediate_reg_0[4564]),.o(intermediate_reg_1[2282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4563]),.i2(intermediate_reg_0[4562]),.o(intermediate_reg_1[2281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4561]),.i2(intermediate_reg_0[4560]),.o(intermediate_reg_1[2280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4559]),.i2(intermediate_reg_0[4558]),.o(intermediate_reg_1[2279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4557]),.i2(intermediate_reg_0[4556]),.o(intermediate_reg_1[2278]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4555]),.i2(intermediate_reg_0[4554]),.o(intermediate_reg_1[2277])); 
mux_module mux_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4553]),.i2(intermediate_reg_0[4552]),.o(intermediate_reg_1[2276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4551]),.i2(intermediate_reg_0[4550]),.o(intermediate_reg_1[2275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4549]),.i2(intermediate_reg_0[4548]),.o(intermediate_reg_1[2274]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4547]),.i2(intermediate_reg_0[4546]),.o(intermediate_reg_1[2273])); 
xor_module xor_module_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4545]),.i2(intermediate_reg_0[4544]),.o(intermediate_reg_1[2272])); 
xor_module xor_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4543]),.i2(intermediate_reg_0[4542]),.o(intermediate_reg_1[2271])); 
xor_module xor_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4541]),.i2(intermediate_reg_0[4540]),.o(intermediate_reg_1[2270])); 
xor_module xor_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4539]),.i2(intermediate_reg_0[4538]),.o(intermediate_reg_1[2269])); 
xor_module xor_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4537]),.i2(intermediate_reg_0[4536]),.o(intermediate_reg_1[2268])); 
mux_module mux_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4535]),.i2(intermediate_reg_0[4534]),.o(intermediate_reg_1[2267]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4533]),.i2(intermediate_reg_0[4532]),.o(intermediate_reg_1[2266]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4531]),.i2(intermediate_reg_0[4530]),.o(intermediate_reg_1[2265])); 
xor_module xor_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4529]),.i2(intermediate_reg_0[4528]),.o(intermediate_reg_1[2264])); 
mux_module mux_module_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4527]),.i2(intermediate_reg_0[4526]),.o(intermediate_reg_1[2263]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4525]),.i2(intermediate_reg_0[4524]),.o(intermediate_reg_1[2262])); 
xor_module xor_module_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4523]),.i2(intermediate_reg_0[4522]),.o(intermediate_reg_1[2261])); 
xor_module xor_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4521]),.i2(intermediate_reg_0[4520]),.o(intermediate_reg_1[2260])); 
mux_module mux_module_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4519]),.i2(intermediate_reg_0[4518]),.o(intermediate_reg_1[2259]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4517]),.i2(intermediate_reg_0[4516]),.o(intermediate_reg_1[2258])); 
mux_module mux_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4515]),.i2(intermediate_reg_0[4514]),.o(intermediate_reg_1[2257]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4513]),.i2(intermediate_reg_0[4512]),.o(intermediate_reg_1[2256])); 
mux_module mux_module_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4511]),.i2(intermediate_reg_0[4510]),.o(intermediate_reg_1[2255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4509]),.i2(intermediate_reg_0[4508]),.o(intermediate_reg_1[2254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4507]),.i2(intermediate_reg_0[4506]),.o(intermediate_reg_1[2253]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4505]),.i2(intermediate_reg_0[4504]),.o(intermediate_reg_1[2252])); 
xor_module xor_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4503]),.i2(intermediate_reg_0[4502]),.o(intermediate_reg_1[2251])); 
xor_module xor_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4501]),.i2(intermediate_reg_0[4500]),.o(intermediate_reg_1[2250])); 
xor_module xor_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4499]),.i2(intermediate_reg_0[4498]),.o(intermediate_reg_1[2249])); 
mux_module mux_module_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4497]),.i2(intermediate_reg_0[4496]),.o(intermediate_reg_1[2248]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4495]),.i2(intermediate_reg_0[4494]),.o(intermediate_reg_1[2247])); 
xor_module xor_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4493]),.i2(intermediate_reg_0[4492]),.o(intermediate_reg_1[2246])); 
mux_module mux_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4491]),.i2(intermediate_reg_0[4490]),.o(intermediate_reg_1[2245]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4489]),.i2(intermediate_reg_0[4488]),.o(intermediate_reg_1[2244])); 
xor_module xor_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4487]),.i2(intermediate_reg_0[4486]),.o(intermediate_reg_1[2243])); 
mux_module mux_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4485]),.i2(intermediate_reg_0[4484]),.o(intermediate_reg_1[2242]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4483]),.i2(intermediate_reg_0[4482]),.o(intermediate_reg_1[2241])); 
mux_module mux_module_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4481]),.i2(intermediate_reg_0[4480]),.o(intermediate_reg_1[2240]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4479]),.i2(intermediate_reg_0[4478]),.o(intermediate_reg_1[2239])); 
xor_module xor_module_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4477]),.i2(intermediate_reg_0[4476]),.o(intermediate_reg_1[2238])); 
xor_module xor_module_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4475]),.i2(intermediate_reg_0[4474]),.o(intermediate_reg_1[2237])); 
mux_module mux_module_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4473]),.i2(intermediate_reg_0[4472]),.o(intermediate_reg_1[2236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4471]),.i2(intermediate_reg_0[4470]),.o(intermediate_reg_1[2235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4469]),.i2(intermediate_reg_0[4468]),.o(intermediate_reg_1[2234]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4467]),.i2(intermediate_reg_0[4466]),.o(intermediate_reg_1[2233])); 
mux_module mux_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4465]),.i2(intermediate_reg_0[4464]),.o(intermediate_reg_1[2232]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4463]),.i2(intermediate_reg_0[4462]),.o(intermediate_reg_1[2231])); 
xor_module xor_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4461]),.i2(intermediate_reg_0[4460]),.o(intermediate_reg_1[2230])); 
xor_module xor_module_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4459]),.i2(intermediate_reg_0[4458]),.o(intermediate_reg_1[2229])); 
xor_module xor_module_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4457]),.i2(intermediate_reg_0[4456]),.o(intermediate_reg_1[2228])); 
mux_module mux_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4455]),.i2(intermediate_reg_0[4454]),.o(intermediate_reg_1[2227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4453]),.i2(intermediate_reg_0[4452]),.o(intermediate_reg_1[2226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4451]),.i2(intermediate_reg_0[4450]),.o(intermediate_reg_1[2225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4449]),.i2(intermediate_reg_0[4448]),.o(intermediate_reg_1[2224])); 
xor_module xor_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4447]),.i2(intermediate_reg_0[4446]),.o(intermediate_reg_1[2223])); 
xor_module xor_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4445]),.i2(intermediate_reg_0[4444]),.o(intermediate_reg_1[2222])); 
mux_module mux_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4443]),.i2(intermediate_reg_0[4442]),.o(intermediate_reg_1[2221]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4441]),.i2(intermediate_reg_0[4440]),.o(intermediate_reg_1[2220]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4439]),.i2(intermediate_reg_0[4438]),.o(intermediate_reg_1[2219])); 
mux_module mux_module_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4437]),.i2(intermediate_reg_0[4436]),.o(intermediate_reg_1[2218]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4435]),.i2(intermediate_reg_0[4434]),.o(intermediate_reg_1[2217]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4433]),.i2(intermediate_reg_0[4432]),.o(intermediate_reg_1[2216])); 
mux_module mux_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4431]),.i2(intermediate_reg_0[4430]),.o(intermediate_reg_1[2215]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4429]),.i2(intermediate_reg_0[4428]),.o(intermediate_reg_1[2214])); 
mux_module mux_module_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4427]),.i2(intermediate_reg_0[4426]),.o(intermediate_reg_1[2213]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4425]),.i2(intermediate_reg_0[4424]),.o(intermediate_reg_1[2212])); 
xor_module xor_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4423]),.i2(intermediate_reg_0[4422]),.o(intermediate_reg_1[2211])); 
mux_module mux_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4421]),.i2(intermediate_reg_0[4420]),.o(intermediate_reg_1[2210]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4419]),.i2(intermediate_reg_0[4418]),.o(intermediate_reg_1[2209]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4417]),.i2(intermediate_reg_0[4416]),.o(intermediate_reg_1[2208]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4415]),.i2(intermediate_reg_0[4414]),.o(intermediate_reg_1[2207])); 
mux_module mux_module_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4413]),.i2(intermediate_reg_0[4412]),.o(intermediate_reg_1[2206]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4411]),.i2(intermediate_reg_0[4410]),.o(intermediate_reg_1[2205])); 
xor_module xor_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4409]),.i2(intermediate_reg_0[4408]),.o(intermediate_reg_1[2204])); 
xor_module xor_module_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4407]),.i2(intermediate_reg_0[4406]),.o(intermediate_reg_1[2203])); 
mux_module mux_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4405]),.i2(intermediate_reg_0[4404]),.o(intermediate_reg_1[2202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4403]),.i2(intermediate_reg_0[4402]),.o(intermediate_reg_1[2201]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4401]),.i2(intermediate_reg_0[4400]),.o(intermediate_reg_1[2200])); 
xor_module xor_module_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4399]),.i2(intermediate_reg_0[4398]),.o(intermediate_reg_1[2199])); 
mux_module mux_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4397]),.i2(intermediate_reg_0[4396]),.o(intermediate_reg_1[2198]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4395]),.i2(intermediate_reg_0[4394]),.o(intermediate_reg_1[2197])); 
xor_module xor_module_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4393]),.i2(intermediate_reg_0[4392]),.o(intermediate_reg_1[2196])); 
xor_module xor_module_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4391]),.i2(intermediate_reg_0[4390]),.o(intermediate_reg_1[2195])); 
xor_module xor_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4389]),.i2(intermediate_reg_0[4388]),.o(intermediate_reg_1[2194])); 
mux_module mux_module_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4387]),.i2(intermediate_reg_0[4386]),.o(intermediate_reg_1[2193]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4385]),.i2(intermediate_reg_0[4384]),.o(intermediate_reg_1[2192])); 
xor_module xor_module_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4383]),.i2(intermediate_reg_0[4382]),.o(intermediate_reg_1[2191])); 
mux_module mux_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4381]),.i2(intermediate_reg_0[4380]),.o(intermediate_reg_1[2190]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4379]),.i2(intermediate_reg_0[4378]),.o(intermediate_reg_1[2189])); 
mux_module mux_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4377]),.i2(intermediate_reg_0[4376]),.o(intermediate_reg_1[2188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4375]),.i2(intermediate_reg_0[4374]),.o(intermediate_reg_1[2187]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4373]),.i2(intermediate_reg_0[4372]),.o(intermediate_reg_1[2186])); 
xor_module xor_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4371]),.i2(intermediate_reg_0[4370]),.o(intermediate_reg_1[2185])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4369]),.i2(intermediate_reg_0[4368]),.o(intermediate_reg_1[2184]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4367]),.i2(intermediate_reg_0[4366]),.o(intermediate_reg_1[2183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4365]),.i2(intermediate_reg_0[4364]),.o(intermediate_reg_1[2182]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4363]),.i2(intermediate_reg_0[4362]),.o(intermediate_reg_1[2181]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4361]),.i2(intermediate_reg_0[4360]),.o(intermediate_reg_1[2180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4359]),.i2(intermediate_reg_0[4358]),.o(intermediate_reg_1[2179]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4357]),.i2(intermediate_reg_0[4356]),.o(intermediate_reg_1[2178])); 
xor_module xor_module_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4355]),.i2(intermediate_reg_0[4354]),.o(intermediate_reg_1[2177])); 
mux_module mux_module_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4353]),.i2(intermediate_reg_0[4352]),.o(intermediate_reg_1[2176]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4351]),.i2(intermediate_reg_0[4350]),.o(intermediate_reg_1[2175])); 
xor_module xor_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4349]),.i2(intermediate_reg_0[4348]),.o(intermediate_reg_1[2174])); 
xor_module xor_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4347]),.i2(intermediate_reg_0[4346]),.o(intermediate_reg_1[2173])); 
mux_module mux_module_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4345]),.i2(intermediate_reg_0[4344]),.o(intermediate_reg_1[2172]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4343]),.i2(intermediate_reg_0[4342]),.o(intermediate_reg_1[2171])); 
mux_module mux_module_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4341]),.i2(intermediate_reg_0[4340]),.o(intermediate_reg_1[2170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4339]),.i2(intermediate_reg_0[4338]),.o(intermediate_reg_1[2169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4337]),.i2(intermediate_reg_0[4336]),.o(intermediate_reg_1[2168]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4335]),.i2(intermediate_reg_0[4334]),.o(intermediate_reg_1[2167])); 
mux_module mux_module_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4333]),.i2(intermediate_reg_0[4332]),.o(intermediate_reg_1[2166]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4331]),.i2(intermediate_reg_0[4330]),.o(intermediate_reg_1[2165])); 
xor_module xor_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4329]),.i2(intermediate_reg_0[4328]),.o(intermediate_reg_1[2164])); 
xor_module xor_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4327]),.i2(intermediate_reg_0[4326]),.o(intermediate_reg_1[2163])); 
xor_module xor_module_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4325]),.i2(intermediate_reg_0[4324]),.o(intermediate_reg_1[2162])); 
mux_module mux_module_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4323]),.i2(intermediate_reg_0[4322]),.o(intermediate_reg_1[2161]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4321]),.i2(intermediate_reg_0[4320]),.o(intermediate_reg_1[2160])); 
xor_module xor_module_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4319]),.i2(intermediate_reg_0[4318]),.o(intermediate_reg_1[2159])); 
mux_module mux_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4317]),.i2(intermediate_reg_0[4316]),.o(intermediate_reg_1[2158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4315]),.i2(intermediate_reg_0[4314]),.o(intermediate_reg_1[2157]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4313]),.i2(intermediate_reg_0[4312]),.o(intermediate_reg_1[2156])); 
xor_module xor_module_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4311]),.i2(intermediate_reg_0[4310]),.o(intermediate_reg_1[2155])); 
xor_module xor_module_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4309]),.i2(intermediate_reg_0[4308]),.o(intermediate_reg_1[2154])); 
xor_module xor_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4307]),.i2(intermediate_reg_0[4306]),.o(intermediate_reg_1[2153])); 
mux_module mux_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4305]),.i2(intermediate_reg_0[4304]),.o(intermediate_reg_1[2152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4303]),.i2(intermediate_reg_0[4302]),.o(intermediate_reg_1[2151]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4301]),.i2(intermediate_reg_0[4300]),.o(intermediate_reg_1[2150])); 
xor_module xor_module_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4299]),.i2(intermediate_reg_0[4298]),.o(intermediate_reg_1[2149])); 
mux_module mux_module_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4297]),.i2(intermediate_reg_0[4296]),.o(intermediate_reg_1[2148]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4295]),.i2(intermediate_reg_0[4294]),.o(intermediate_reg_1[2147])); 
mux_module mux_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4293]),.i2(intermediate_reg_0[4292]),.o(intermediate_reg_1[2146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4291]),.i2(intermediate_reg_0[4290]),.o(intermediate_reg_1[2145]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4289]),.i2(intermediate_reg_0[4288]),.o(intermediate_reg_1[2144])); 
mux_module mux_module_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4287]),.i2(intermediate_reg_0[4286]),.o(intermediate_reg_1[2143]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4285]),.i2(intermediate_reg_0[4284]),.o(intermediate_reg_1[2142])); 
mux_module mux_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4283]),.i2(intermediate_reg_0[4282]),.o(intermediate_reg_1[2141]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4281]),.i2(intermediate_reg_0[4280]),.o(intermediate_reg_1[2140])); 
mux_module mux_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4279]),.i2(intermediate_reg_0[4278]),.o(intermediate_reg_1[2139]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4277]),.i2(intermediate_reg_0[4276]),.o(intermediate_reg_1[2138]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4275]),.i2(intermediate_reg_0[4274]),.o(intermediate_reg_1[2137])); 
xor_module xor_module_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4273]),.i2(intermediate_reg_0[4272]),.o(intermediate_reg_1[2136])); 
mux_module mux_module_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4271]),.i2(intermediate_reg_0[4270]),.o(intermediate_reg_1[2135]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4269]),.i2(intermediate_reg_0[4268]),.o(intermediate_reg_1[2134])); 
xor_module xor_module_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4267]),.i2(intermediate_reg_0[4266]),.o(intermediate_reg_1[2133])); 
mux_module mux_module_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4265]),.i2(intermediate_reg_0[4264]),.o(intermediate_reg_1[2132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4263]),.i2(intermediate_reg_0[4262]),.o(intermediate_reg_1[2131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4261]),.i2(intermediate_reg_0[4260]),.o(intermediate_reg_1[2130]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4259]),.i2(intermediate_reg_0[4258]),.o(intermediate_reg_1[2129]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4257]),.i2(intermediate_reg_0[4256]),.o(intermediate_reg_1[2128])); 
xor_module xor_module_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4255]),.i2(intermediate_reg_0[4254]),.o(intermediate_reg_1[2127])); 
mux_module mux_module_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4253]),.i2(intermediate_reg_0[4252]),.o(intermediate_reg_1[2126]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4251]),.i2(intermediate_reg_0[4250]),.o(intermediate_reg_1[2125]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4249]),.i2(intermediate_reg_0[4248]),.o(intermediate_reg_1[2124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4247]),.i2(intermediate_reg_0[4246]),.o(intermediate_reg_1[2123]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4245]),.i2(intermediate_reg_0[4244]),.o(intermediate_reg_1[2122])); 
xor_module xor_module_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4243]),.i2(intermediate_reg_0[4242]),.o(intermediate_reg_1[2121])); 
mux_module mux_module_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4241]),.i2(intermediate_reg_0[4240]),.o(intermediate_reg_1[2120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4239]),.i2(intermediate_reg_0[4238]),.o(intermediate_reg_1[2119]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4237]),.i2(intermediate_reg_0[4236]),.o(intermediate_reg_1[2118]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4235]),.i2(intermediate_reg_0[4234]),.o(intermediate_reg_1[2117])); 
xor_module xor_module_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4233]),.i2(intermediate_reg_0[4232]),.o(intermediate_reg_1[2116])); 
xor_module xor_module_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4231]),.i2(intermediate_reg_0[4230]),.o(intermediate_reg_1[2115])); 
xor_module xor_module_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4229]),.i2(intermediate_reg_0[4228]),.o(intermediate_reg_1[2114])); 
mux_module mux_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4227]),.i2(intermediate_reg_0[4226]),.o(intermediate_reg_1[2113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4225]),.i2(intermediate_reg_0[4224]),.o(intermediate_reg_1[2112]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4223]),.i2(intermediate_reg_0[4222]),.o(intermediate_reg_1[2111])); 
mux_module mux_module_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4221]),.i2(intermediate_reg_0[4220]),.o(intermediate_reg_1[2110]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4219]),.i2(intermediate_reg_0[4218]),.o(intermediate_reg_1[2109]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4217]),.i2(intermediate_reg_0[4216]),.o(intermediate_reg_1[2108])); 
xor_module xor_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4215]),.i2(intermediate_reg_0[4214]),.o(intermediate_reg_1[2107])); 
mux_module mux_module_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4213]),.i2(intermediate_reg_0[4212]),.o(intermediate_reg_1[2106]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4211]),.i2(intermediate_reg_0[4210]),.o(intermediate_reg_1[2105]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4209]),.i2(intermediate_reg_0[4208]),.o(intermediate_reg_1[2104]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4207]),.i2(intermediate_reg_0[4206]),.o(intermediate_reg_1[2103])); 
mux_module mux_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4205]),.i2(intermediate_reg_0[4204]),.o(intermediate_reg_1[2102]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4203]),.i2(intermediate_reg_0[4202]),.o(intermediate_reg_1[2101])); 
mux_module mux_module_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4201]),.i2(intermediate_reg_0[4200]),.o(intermediate_reg_1[2100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4199]),.i2(intermediate_reg_0[4198]),.o(intermediate_reg_1[2099]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4197]),.i2(intermediate_reg_0[4196]),.o(intermediate_reg_1[2098])); 
mux_module mux_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4195]),.i2(intermediate_reg_0[4194]),.o(intermediate_reg_1[2097]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4193]),.i2(intermediate_reg_0[4192]),.o(intermediate_reg_1[2096])); 
mux_module mux_module_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4191]),.i2(intermediate_reg_0[4190]),.o(intermediate_reg_1[2095]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4189]),.i2(intermediate_reg_0[4188]),.o(intermediate_reg_1[2094]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4187]),.i2(intermediate_reg_0[4186]),.o(intermediate_reg_1[2093]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4185]),.i2(intermediate_reg_0[4184]),.o(intermediate_reg_1[2092])); 
mux_module mux_module_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4183]),.i2(intermediate_reg_0[4182]),.o(intermediate_reg_1[2091]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4181]),.i2(intermediate_reg_0[4180]),.o(intermediate_reg_1[2090]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4179]),.i2(intermediate_reg_0[4178]),.o(intermediate_reg_1[2089])); 
mux_module mux_module_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4177]),.i2(intermediate_reg_0[4176]),.o(intermediate_reg_1[2088]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4175]),.i2(intermediate_reg_0[4174]),.o(intermediate_reg_1[2087]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4173]),.i2(intermediate_reg_0[4172]),.o(intermediate_reg_1[2086]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4171]),.i2(intermediate_reg_0[4170]),.o(intermediate_reg_1[2085]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4169]),.i2(intermediate_reg_0[4168]),.o(intermediate_reg_1[2084]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4167]),.i2(intermediate_reg_0[4166]),.o(intermediate_reg_1[2083]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4165]),.i2(intermediate_reg_0[4164]),.o(intermediate_reg_1[2082])); 
mux_module mux_module_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4163]),.i2(intermediate_reg_0[4162]),.o(intermediate_reg_1[2081]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4161]),.i2(intermediate_reg_0[4160]),.o(intermediate_reg_1[2080])); 
xor_module xor_module_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4159]),.i2(intermediate_reg_0[4158]),.o(intermediate_reg_1[2079])); 
mux_module mux_module_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4157]),.i2(intermediate_reg_0[4156]),.o(intermediate_reg_1[2078]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4155]),.i2(intermediate_reg_0[4154]),.o(intermediate_reg_1[2077]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4153]),.i2(intermediate_reg_0[4152]),.o(intermediate_reg_1[2076])); 
xor_module xor_module_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4151]),.i2(intermediate_reg_0[4150]),.o(intermediate_reg_1[2075])); 
mux_module mux_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4149]),.i2(intermediate_reg_0[4148]),.o(intermediate_reg_1[2074]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4147]),.i2(intermediate_reg_0[4146]),.o(intermediate_reg_1[2073]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4145]),.i2(intermediate_reg_0[4144]),.o(intermediate_reg_1[2072])); 
xor_module xor_module_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4143]),.i2(intermediate_reg_0[4142]),.o(intermediate_reg_1[2071])); 
mux_module mux_module_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4141]),.i2(intermediate_reg_0[4140]),.o(intermediate_reg_1[2070]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4139]),.i2(intermediate_reg_0[4138]),.o(intermediate_reg_1[2069])); 
xor_module xor_module_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4137]),.i2(intermediate_reg_0[4136]),.o(intermediate_reg_1[2068])); 
xor_module xor_module_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4135]),.i2(intermediate_reg_0[4134]),.o(intermediate_reg_1[2067])); 
xor_module xor_module_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4133]),.i2(intermediate_reg_0[4132]),.o(intermediate_reg_1[2066])); 
xor_module xor_module_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4131]),.i2(intermediate_reg_0[4130]),.o(intermediate_reg_1[2065])); 
mux_module mux_module_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4129]),.i2(intermediate_reg_0[4128]),.o(intermediate_reg_1[2064]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4127]),.i2(intermediate_reg_0[4126]),.o(intermediate_reg_1[2063])); 
xor_module xor_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4125]),.i2(intermediate_reg_0[4124]),.o(intermediate_reg_1[2062])); 
xor_module xor_module_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4123]),.i2(intermediate_reg_0[4122]),.o(intermediate_reg_1[2061])); 
mux_module mux_module_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4121]),.i2(intermediate_reg_0[4120]),.o(intermediate_reg_1[2060]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4119]),.i2(intermediate_reg_0[4118]),.o(intermediate_reg_1[2059]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4117]),.i2(intermediate_reg_0[4116]),.o(intermediate_reg_1[2058])); 
xor_module xor_module_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4115]),.i2(intermediate_reg_0[4114]),.o(intermediate_reg_1[2057])); 
mux_module mux_module_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4113]),.i2(intermediate_reg_0[4112]),.o(intermediate_reg_1[2056]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4111]),.i2(intermediate_reg_0[4110]),.o(intermediate_reg_1[2055])); 
mux_module mux_module_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4109]),.i2(intermediate_reg_0[4108]),.o(intermediate_reg_1[2054]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4107]),.i2(intermediate_reg_0[4106]),.o(intermediate_reg_1[2053]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4105]),.i2(intermediate_reg_0[4104]),.o(intermediate_reg_1[2052])); 
mux_module mux_module_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4103]),.i2(intermediate_reg_0[4102]),.o(intermediate_reg_1[2051]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4101]),.i2(intermediate_reg_0[4100]),.o(intermediate_reg_1[2050]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4099]),.i2(intermediate_reg_0[4098]),.o(intermediate_reg_1[2049])); 
xor_module xor_module_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4097]),.i2(intermediate_reg_0[4096]),.o(intermediate_reg_1[2048])); 
xor_module xor_module_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4095]),.i2(intermediate_reg_0[4094]),.o(intermediate_reg_1[2047])); 
xor_module xor_module_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4093]),.i2(intermediate_reg_0[4092]),.o(intermediate_reg_1[2046])); 
mux_module mux_module_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4091]),.i2(intermediate_reg_0[4090]),.o(intermediate_reg_1[2045]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4089]),.i2(intermediate_reg_0[4088]),.o(intermediate_reg_1[2044])); 
mux_module mux_module_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4087]),.i2(intermediate_reg_0[4086]),.o(intermediate_reg_1[2043]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4085]),.i2(intermediate_reg_0[4084]),.o(intermediate_reg_1[2042]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4083]),.i2(intermediate_reg_0[4082]),.o(intermediate_reg_1[2041])); 
xor_module xor_module_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4081]),.i2(intermediate_reg_0[4080]),.o(intermediate_reg_1[2040])); 
xor_module xor_module_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4079]),.i2(intermediate_reg_0[4078]),.o(intermediate_reg_1[2039])); 
mux_module mux_module_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4077]),.i2(intermediate_reg_0[4076]),.o(intermediate_reg_1[2038]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4075]),.i2(intermediate_reg_0[4074]),.o(intermediate_reg_1[2037]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4073]),.i2(intermediate_reg_0[4072]),.o(intermediate_reg_1[2036]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4071]),.i2(intermediate_reg_0[4070]),.o(intermediate_reg_1[2035]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4069]),.i2(intermediate_reg_0[4068]),.o(intermediate_reg_1[2034])); 
mux_module mux_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4067]),.i2(intermediate_reg_0[4066]),.o(intermediate_reg_1[2033]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4065]),.i2(intermediate_reg_0[4064]),.o(intermediate_reg_1[2032]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4063]),.i2(intermediate_reg_0[4062]),.o(intermediate_reg_1[2031])); 
mux_module mux_module_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4061]),.i2(intermediate_reg_0[4060]),.o(intermediate_reg_1[2030]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4059]),.i2(intermediate_reg_0[4058]),.o(intermediate_reg_1[2029]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4057]),.i2(intermediate_reg_0[4056]),.o(intermediate_reg_1[2028])); 
mux_module mux_module_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4055]),.i2(intermediate_reg_0[4054]),.o(intermediate_reg_1[2027]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4053]),.i2(intermediate_reg_0[4052]),.o(intermediate_reg_1[2026]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4051]),.i2(intermediate_reg_0[4050]),.o(intermediate_reg_1[2025])); 
mux_module mux_module_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4049]),.i2(intermediate_reg_0[4048]),.o(intermediate_reg_1[2024]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4047]),.i2(intermediate_reg_0[4046]),.o(intermediate_reg_1[2023])); 
mux_module mux_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4045]),.i2(intermediate_reg_0[4044]),.o(intermediate_reg_1[2022]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4043]),.i2(intermediate_reg_0[4042]),.o(intermediate_reg_1[2021]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4041]),.i2(intermediate_reg_0[4040]),.o(intermediate_reg_1[2020]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4039]),.i2(intermediate_reg_0[4038]),.o(intermediate_reg_1[2019]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4037]),.i2(intermediate_reg_0[4036]),.o(intermediate_reg_1[2018])); 
xor_module xor_module_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4035]),.i2(intermediate_reg_0[4034]),.o(intermediate_reg_1[2017])); 
xor_module xor_module_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4033]),.i2(intermediate_reg_0[4032]),.o(intermediate_reg_1[2016])); 
mux_module mux_module_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4031]),.i2(intermediate_reg_0[4030]),.o(intermediate_reg_1[2015]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4029]),.i2(intermediate_reg_0[4028]),.o(intermediate_reg_1[2014]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4027]),.i2(intermediate_reg_0[4026]),.o(intermediate_reg_1[2013]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4025]),.i2(intermediate_reg_0[4024]),.o(intermediate_reg_1[2012])); 
mux_module mux_module_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4023]),.i2(intermediate_reg_0[4022]),.o(intermediate_reg_1[2011]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4021]),.i2(intermediate_reg_0[4020]),.o(intermediate_reg_1[2010])); 
xor_module xor_module_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4019]),.i2(intermediate_reg_0[4018]),.o(intermediate_reg_1[2009])); 
xor_module xor_module_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4017]),.i2(intermediate_reg_0[4016]),.o(intermediate_reg_1[2008])); 
xor_module xor_module_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4015]),.i2(intermediate_reg_0[4014]),.o(intermediate_reg_1[2007])); 
mux_module mux_module_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4013]),.i2(intermediate_reg_0[4012]),.o(intermediate_reg_1[2006]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4011]),.i2(intermediate_reg_0[4010]),.o(intermediate_reg_1[2005]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4009]),.i2(intermediate_reg_0[4008]),.o(intermediate_reg_1[2004]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4007]),.i2(intermediate_reg_0[4006]),.o(intermediate_reg_1[2003]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4005]),.i2(intermediate_reg_0[4004]),.o(intermediate_reg_1[2002]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4003]),.i2(intermediate_reg_0[4002]),.o(intermediate_reg_1[2001])); 
mux_module mux_module_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4001]),.i2(intermediate_reg_0[4000]),.o(intermediate_reg_1[2000]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3999]),.i2(intermediate_reg_0[3998]),.o(intermediate_reg_1[1999])); 
mux_module mux_module_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3997]),.i2(intermediate_reg_0[3996]),.o(intermediate_reg_1[1998]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3995]),.i2(intermediate_reg_0[3994]),.o(intermediate_reg_1[1997])); 
xor_module xor_module_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3993]),.i2(intermediate_reg_0[3992]),.o(intermediate_reg_1[1996])); 
mux_module mux_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3991]),.i2(intermediate_reg_0[3990]),.o(intermediate_reg_1[1995]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3989]),.i2(intermediate_reg_0[3988]),.o(intermediate_reg_1[1994])); 
xor_module xor_module_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3987]),.i2(intermediate_reg_0[3986]),.o(intermediate_reg_1[1993])); 
xor_module xor_module_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3985]),.i2(intermediate_reg_0[3984]),.o(intermediate_reg_1[1992])); 
mux_module mux_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3983]),.i2(intermediate_reg_0[3982]),.o(intermediate_reg_1[1991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3981]),.i2(intermediate_reg_0[3980]),.o(intermediate_reg_1[1990]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3979]),.i2(intermediate_reg_0[3978]),.o(intermediate_reg_1[1989])); 
mux_module mux_module_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3977]),.i2(intermediate_reg_0[3976]),.o(intermediate_reg_1[1988]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3975]),.i2(intermediate_reg_0[3974]),.o(intermediate_reg_1[1987]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3973]),.i2(intermediate_reg_0[3972]),.o(intermediate_reg_1[1986])); 
xor_module xor_module_inst_1_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3971]),.i2(intermediate_reg_0[3970]),.o(intermediate_reg_1[1985])); 
xor_module xor_module_inst_1_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3969]),.i2(intermediate_reg_0[3968]),.o(intermediate_reg_1[1984])); 
xor_module xor_module_inst_1_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3967]),.i2(intermediate_reg_0[3966]),.o(intermediate_reg_1[1983])); 
xor_module xor_module_inst_1_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3965]),.i2(intermediate_reg_0[3964]),.o(intermediate_reg_1[1982])); 
xor_module xor_module_inst_1_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3963]),.i2(intermediate_reg_0[3962]),.o(intermediate_reg_1[1981])); 
xor_module xor_module_inst_1_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3961]),.i2(intermediate_reg_0[3960]),.o(intermediate_reg_1[1980])); 
mux_module mux_module_inst_1_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3959]),.i2(intermediate_reg_0[3958]),.o(intermediate_reg_1[1979]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3957]),.i2(intermediate_reg_0[3956]),.o(intermediate_reg_1[1978]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3955]),.i2(intermediate_reg_0[3954]),.o(intermediate_reg_1[1977]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3953]),.i2(intermediate_reg_0[3952]),.o(intermediate_reg_1[1976]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3951]),.i2(intermediate_reg_0[3950]),.o(intermediate_reg_1[1975])); 
xor_module xor_module_inst_1_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3949]),.i2(intermediate_reg_0[3948]),.o(intermediate_reg_1[1974])); 
mux_module mux_module_inst_1_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3947]),.i2(intermediate_reg_0[3946]),.o(intermediate_reg_1[1973]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3945]),.i2(intermediate_reg_0[3944]),.o(intermediate_reg_1[1972]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3943]),.i2(intermediate_reg_0[3942]),.o(intermediate_reg_1[1971]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3941]),.i2(intermediate_reg_0[3940]),.o(intermediate_reg_1[1970])); 
xor_module xor_module_inst_1_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3939]),.i2(intermediate_reg_0[3938]),.o(intermediate_reg_1[1969])); 
xor_module xor_module_inst_1_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3937]),.i2(intermediate_reg_0[3936]),.o(intermediate_reg_1[1968])); 
mux_module mux_module_inst_1_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3935]),.i2(intermediate_reg_0[3934]),.o(intermediate_reg_1[1967]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3933]),.i2(intermediate_reg_0[3932]),.o(intermediate_reg_1[1966]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3931]),.i2(intermediate_reg_0[3930]),.o(intermediate_reg_1[1965]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3929]),.i2(intermediate_reg_0[3928]),.o(intermediate_reg_1[1964])); 
mux_module mux_module_inst_1_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3927]),.i2(intermediate_reg_0[3926]),.o(intermediate_reg_1[1963]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3925]),.i2(intermediate_reg_0[3924]),.o(intermediate_reg_1[1962])); 
xor_module xor_module_inst_1_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3923]),.i2(intermediate_reg_0[3922]),.o(intermediate_reg_1[1961])); 
mux_module mux_module_inst_1_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3921]),.i2(intermediate_reg_0[3920]),.o(intermediate_reg_1[1960]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3919]),.i2(intermediate_reg_0[3918]),.o(intermediate_reg_1[1959]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3917]),.i2(intermediate_reg_0[3916]),.o(intermediate_reg_1[1958])); 
xor_module xor_module_inst_1_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3915]),.i2(intermediate_reg_0[3914]),.o(intermediate_reg_1[1957])); 
xor_module xor_module_inst_1_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3913]),.i2(intermediate_reg_0[3912]),.o(intermediate_reg_1[1956])); 
mux_module mux_module_inst_1_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3911]),.i2(intermediate_reg_0[3910]),.o(intermediate_reg_1[1955]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3909]),.i2(intermediate_reg_0[3908]),.o(intermediate_reg_1[1954])); 
mux_module mux_module_inst_1_1344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3907]),.i2(intermediate_reg_0[3906]),.o(intermediate_reg_1[1953]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3905]),.i2(intermediate_reg_0[3904]),.o(intermediate_reg_1[1952]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3903]),.i2(intermediate_reg_0[3902]),.o(intermediate_reg_1[1951]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3901]),.i2(intermediate_reg_0[3900]),.o(intermediate_reg_1[1950])); 
xor_module xor_module_inst_1_1348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3899]),.i2(intermediate_reg_0[3898]),.o(intermediate_reg_1[1949])); 
mux_module mux_module_inst_1_1349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3897]),.i2(intermediate_reg_0[3896]),.o(intermediate_reg_1[1948]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3895]),.i2(intermediate_reg_0[3894]),.o(intermediate_reg_1[1947]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3893]),.i2(intermediate_reg_0[3892]),.o(intermediate_reg_1[1946]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3891]),.i2(intermediate_reg_0[3890]),.o(intermediate_reg_1[1945])); 
mux_module mux_module_inst_1_1353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3889]),.i2(intermediate_reg_0[3888]),.o(intermediate_reg_1[1944]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3887]),.i2(intermediate_reg_0[3886]),.o(intermediate_reg_1[1943])); 
mux_module mux_module_inst_1_1355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3885]),.i2(intermediate_reg_0[3884]),.o(intermediate_reg_1[1942]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3883]),.i2(intermediate_reg_0[3882]),.o(intermediate_reg_1[1941])); 
xor_module xor_module_inst_1_1357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3881]),.i2(intermediate_reg_0[3880]),.o(intermediate_reg_1[1940])); 
xor_module xor_module_inst_1_1358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3879]),.i2(intermediate_reg_0[3878]),.o(intermediate_reg_1[1939])); 
xor_module xor_module_inst_1_1359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3877]),.i2(intermediate_reg_0[3876]),.o(intermediate_reg_1[1938])); 
xor_module xor_module_inst_1_1360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3875]),.i2(intermediate_reg_0[3874]),.o(intermediate_reg_1[1937])); 
xor_module xor_module_inst_1_1361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3873]),.i2(intermediate_reg_0[3872]),.o(intermediate_reg_1[1936])); 
xor_module xor_module_inst_1_1362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3871]),.i2(intermediate_reg_0[3870]),.o(intermediate_reg_1[1935])); 
xor_module xor_module_inst_1_1363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3869]),.i2(intermediate_reg_0[3868]),.o(intermediate_reg_1[1934])); 
xor_module xor_module_inst_1_1364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3867]),.i2(intermediate_reg_0[3866]),.o(intermediate_reg_1[1933])); 
mux_module mux_module_inst_1_1365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3865]),.i2(intermediate_reg_0[3864]),.o(intermediate_reg_1[1932]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3863]),.i2(intermediate_reg_0[3862]),.o(intermediate_reg_1[1931]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3861]),.i2(intermediate_reg_0[3860]),.o(intermediate_reg_1[1930]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3859]),.i2(intermediate_reg_0[3858]),.o(intermediate_reg_1[1929]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3857]),.i2(intermediate_reg_0[3856]),.o(intermediate_reg_1[1928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3855]),.i2(intermediate_reg_0[3854]),.o(intermediate_reg_1[1927]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3853]),.i2(intermediate_reg_0[3852]),.o(intermediate_reg_1[1926]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3851]),.i2(intermediate_reg_0[3850]),.o(intermediate_reg_1[1925]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3849]),.i2(intermediate_reg_0[3848]),.o(intermediate_reg_1[1924]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3847]),.i2(intermediate_reg_0[3846]),.o(intermediate_reg_1[1923])); 
mux_module mux_module_inst_1_1375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3845]),.i2(intermediate_reg_0[3844]),.o(intermediate_reg_1[1922]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3843]),.i2(intermediate_reg_0[3842]),.o(intermediate_reg_1[1921]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3841]),.i2(intermediate_reg_0[3840]),.o(intermediate_reg_1[1920]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3839]),.i2(intermediate_reg_0[3838]),.o(intermediate_reg_1[1919]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3837]),.i2(intermediate_reg_0[3836]),.o(intermediate_reg_1[1918]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3835]),.i2(intermediate_reg_0[3834]),.o(intermediate_reg_1[1917])); 
xor_module xor_module_inst_1_1381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3833]),.i2(intermediate_reg_0[3832]),.o(intermediate_reg_1[1916])); 
mux_module mux_module_inst_1_1382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3831]),.i2(intermediate_reg_0[3830]),.o(intermediate_reg_1[1915]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3829]),.i2(intermediate_reg_0[3828]),.o(intermediate_reg_1[1914]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3827]),.i2(intermediate_reg_0[3826]),.o(intermediate_reg_1[1913]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3825]),.i2(intermediate_reg_0[3824]),.o(intermediate_reg_1[1912])); 
xor_module xor_module_inst_1_1386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3823]),.i2(intermediate_reg_0[3822]),.o(intermediate_reg_1[1911])); 
xor_module xor_module_inst_1_1387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3821]),.i2(intermediate_reg_0[3820]),.o(intermediate_reg_1[1910])); 
mux_module mux_module_inst_1_1388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3819]),.i2(intermediate_reg_0[3818]),.o(intermediate_reg_1[1909]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3817]),.i2(intermediate_reg_0[3816]),.o(intermediate_reg_1[1908]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3815]),.i2(intermediate_reg_0[3814]),.o(intermediate_reg_1[1907]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3813]),.i2(intermediate_reg_0[3812]),.o(intermediate_reg_1[1906]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3811]),.i2(intermediate_reg_0[3810]),.o(intermediate_reg_1[1905])); 
mux_module mux_module_inst_1_1393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3809]),.i2(intermediate_reg_0[3808]),.o(intermediate_reg_1[1904]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3807]),.i2(intermediate_reg_0[3806]),.o(intermediate_reg_1[1903])); 
xor_module xor_module_inst_1_1395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3805]),.i2(intermediate_reg_0[3804]),.o(intermediate_reg_1[1902])); 
xor_module xor_module_inst_1_1396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3803]),.i2(intermediate_reg_0[3802]),.o(intermediate_reg_1[1901])); 
xor_module xor_module_inst_1_1397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3801]),.i2(intermediate_reg_0[3800]),.o(intermediate_reg_1[1900])); 
xor_module xor_module_inst_1_1398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3799]),.i2(intermediate_reg_0[3798]),.o(intermediate_reg_1[1899])); 
xor_module xor_module_inst_1_1399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3797]),.i2(intermediate_reg_0[3796]),.o(intermediate_reg_1[1898])); 
xor_module xor_module_inst_1_1400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3795]),.i2(intermediate_reg_0[3794]),.o(intermediate_reg_1[1897])); 
xor_module xor_module_inst_1_1401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3793]),.i2(intermediate_reg_0[3792]),.o(intermediate_reg_1[1896])); 
mux_module mux_module_inst_1_1402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3791]),.i2(intermediate_reg_0[3790]),.o(intermediate_reg_1[1895]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3789]),.i2(intermediate_reg_0[3788]),.o(intermediate_reg_1[1894])); 
mux_module mux_module_inst_1_1404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3787]),.i2(intermediate_reg_0[3786]),.o(intermediate_reg_1[1893]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3785]),.i2(intermediate_reg_0[3784]),.o(intermediate_reg_1[1892])); 
mux_module mux_module_inst_1_1406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3783]),.i2(intermediate_reg_0[3782]),.o(intermediate_reg_1[1891]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3781]),.i2(intermediate_reg_0[3780]),.o(intermediate_reg_1[1890])); 
xor_module xor_module_inst_1_1408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3779]),.i2(intermediate_reg_0[3778]),.o(intermediate_reg_1[1889])); 
xor_module xor_module_inst_1_1409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3777]),.i2(intermediate_reg_0[3776]),.o(intermediate_reg_1[1888])); 
mux_module mux_module_inst_1_1410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3775]),.i2(intermediate_reg_0[3774]),.o(intermediate_reg_1[1887]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3773]),.i2(intermediate_reg_0[3772]),.o(intermediate_reg_1[1886])); 
xor_module xor_module_inst_1_1412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3771]),.i2(intermediate_reg_0[3770]),.o(intermediate_reg_1[1885])); 
mux_module mux_module_inst_1_1413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3769]),.i2(intermediate_reg_0[3768]),.o(intermediate_reg_1[1884]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3767]),.i2(intermediate_reg_0[3766]),.o(intermediate_reg_1[1883]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3765]),.i2(intermediate_reg_0[3764]),.o(intermediate_reg_1[1882])); 
mux_module mux_module_inst_1_1416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3763]),.i2(intermediate_reg_0[3762]),.o(intermediate_reg_1[1881]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3761]),.i2(intermediate_reg_0[3760]),.o(intermediate_reg_1[1880]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3759]),.i2(intermediate_reg_0[3758]),.o(intermediate_reg_1[1879]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3757]),.i2(intermediate_reg_0[3756]),.o(intermediate_reg_1[1878])); 
mux_module mux_module_inst_1_1420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3755]),.i2(intermediate_reg_0[3754]),.o(intermediate_reg_1[1877]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3753]),.i2(intermediate_reg_0[3752]),.o(intermediate_reg_1[1876]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3751]),.i2(intermediate_reg_0[3750]),.o(intermediate_reg_1[1875])); 
xor_module xor_module_inst_1_1423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3749]),.i2(intermediate_reg_0[3748]),.o(intermediate_reg_1[1874])); 
mux_module mux_module_inst_1_1424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3747]),.i2(intermediate_reg_0[3746]),.o(intermediate_reg_1[1873]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3745]),.i2(intermediate_reg_0[3744]),.o(intermediate_reg_1[1872]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3743]),.i2(intermediate_reg_0[3742]),.o(intermediate_reg_1[1871]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3741]),.i2(intermediate_reg_0[3740]),.o(intermediate_reg_1[1870]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3739]),.i2(intermediate_reg_0[3738]),.o(intermediate_reg_1[1869]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3737]),.i2(intermediate_reg_0[3736]),.o(intermediate_reg_1[1868])); 
mux_module mux_module_inst_1_1430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3735]),.i2(intermediate_reg_0[3734]),.o(intermediate_reg_1[1867]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3733]),.i2(intermediate_reg_0[3732]),.o(intermediate_reg_1[1866])); 
mux_module mux_module_inst_1_1432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3731]),.i2(intermediate_reg_0[3730]),.o(intermediate_reg_1[1865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3729]),.i2(intermediate_reg_0[3728]),.o(intermediate_reg_1[1864]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3727]),.i2(intermediate_reg_0[3726]),.o(intermediate_reg_1[1863])); 
xor_module xor_module_inst_1_1435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3725]),.i2(intermediate_reg_0[3724]),.o(intermediate_reg_1[1862])); 
mux_module mux_module_inst_1_1436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3723]),.i2(intermediate_reg_0[3722]),.o(intermediate_reg_1[1861]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3721]),.i2(intermediate_reg_0[3720]),.o(intermediate_reg_1[1860])); 
xor_module xor_module_inst_1_1438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3719]),.i2(intermediate_reg_0[3718]),.o(intermediate_reg_1[1859])); 
xor_module xor_module_inst_1_1439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3717]),.i2(intermediate_reg_0[3716]),.o(intermediate_reg_1[1858])); 
mux_module mux_module_inst_1_1440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3715]),.i2(intermediate_reg_0[3714]),.o(intermediate_reg_1[1857]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3713]),.i2(intermediate_reg_0[3712]),.o(intermediate_reg_1[1856])); 
xor_module xor_module_inst_1_1442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3711]),.i2(intermediate_reg_0[3710]),.o(intermediate_reg_1[1855])); 
xor_module xor_module_inst_1_1443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3709]),.i2(intermediate_reg_0[3708]),.o(intermediate_reg_1[1854])); 
mux_module mux_module_inst_1_1444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3707]),.i2(intermediate_reg_0[3706]),.o(intermediate_reg_1[1853]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3705]),.i2(intermediate_reg_0[3704]),.o(intermediate_reg_1[1852])); 
xor_module xor_module_inst_1_1446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3703]),.i2(intermediate_reg_0[3702]),.o(intermediate_reg_1[1851])); 
mux_module mux_module_inst_1_1447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3701]),.i2(intermediate_reg_0[3700]),.o(intermediate_reg_1[1850]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3699]),.i2(intermediate_reg_0[3698]),.o(intermediate_reg_1[1849])); 
mux_module mux_module_inst_1_1449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3697]),.i2(intermediate_reg_0[3696]),.o(intermediate_reg_1[1848]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3695]),.i2(intermediate_reg_0[3694]),.o(intermediate_reg_1[1847]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3693]),.i2(intermediate_reg_0[3692]),.o(intermediate_reg_1[1846]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3691]),.i2(intermediate_reg_0[3690]),.o(intermediate_reg_1[1845]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3689]),.i2(intermediate_reg_0[3688]),.o(intermediate_reg_1[1844])); 
xor_module xor_module_inst_1_1454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3687]),.i2(intermediate_reg_0[3686]),.o(intermediate_reg_1[1843])); 
mux_module mux_module_inst_1_1455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3685]),.i2(intermediate_reg_0[3684]),.o(intermediate_reg_1[1842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3683]),.i2(intermediate_reg_0[3682]),.o(intermediate_reg_1[1841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3681]),.i2(intermediate_reg_0[3680]),.o(intermediate_reg_1[1840]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3679]),.i2(intermediate_reg_0[3678]),.o(intermediate_reg_1[1839]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3677]),.i2(intermediate_reg_0[3676]),.o(intermediate_reg_1[1838]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3675]),.i2(intermediate_reg_0[3674]),.o(intermediate_reg_1[1837]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3673]),.i2(intermediate_reg_0[3672]),.o(intermediate_reg_1[1836])); 
xor_module xor_module_inst_1_1462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3671]),.i2(intermediate_reg_0[3670]),.o(intermediate_reg_1[1835])); 
xor_module xor_module_inst_1_1463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3669]),.i2(intermediate_reg_0[3668]),.o(intermediate_reg_1[1834])); 
mux_module mux_module_inst_1_1464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3667]),.i2(intermediate_reg_0[3666]),.o(intermediate_reg_1[1833]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3665]),.i2(intermediate_reg_0[3664]),.o(intermediate_reg_1[1832]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3663]),.i2(intermediate_reg_0[3662]),.o(intermediate_reg_1[1831])); 
mux_module mux_module_inst_1_1467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3661]),.i2(intermediate_reg_0[3660]),.o(intermediate_reg_1[1830]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3659]),.i2(intermediate_reg_0[3658]),.o(intermediate_reg_1[1829])); 
mux_module mux_module_inst_1_1469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3657]),.i2(intermediate_reg_0[3656]),.o(intermediate_reg_1[1828]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3655]),.i2(intermediate_reg_0[3654]),.o(intermediate_reg_1[1827]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3653]),.i2(intermediate_reg_0[3652]),.o(intermediate_reg_1[1826])); 
xor_module xor_module_inst_1_1472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3651]),.i2(intermediate_reg_0[3650]),.o(intermediate_reg_1[1825])); 
mux_module mux_module_inst_1_1473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3649]),.i2(intermediate_reg_0[3648]),.o(intermediate_reg_1[1824]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3647]),.i2(intermediate_reg_0[3646]),.o(intermediate_reg_1[1823])); 
xor_module xor_module_inst_1_1475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3645]),.i2(intermediate_reg_0[3644]),.o(intermediate_reg_1[1822])); 
mux_module mux_module_inst_1_1476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3643]),.i2(intermediate_reg_0[3642]),.o(intermediate_reg_1[1821]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3641]),.i2(intermediate_reg_0[3640]),.o(intermediate_reg_1[1820])); 
mux_module mux_module_inst_1_1478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3639]),.i2(intermediate_reg_0[3638]),.o(intermediate_reg_1[1819]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3637]),.i2(intermediate_reg_0[3636]),.o(intermediate_reg_1[1818]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3635]),.i2(intermediate_reg_0[3634]),.o(intermediate_reg_1[1817]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3633]),.i2(intermediate_reg_0[3632]),.o(intermediate_reg_1[1816]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3631]),.i2(intermediate_reg_0[3630]),.o(intermediate_reg_1[1815]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3629]),.i2(intermediate_reg_0[3628]),.o(intermediate_reg_1[1814]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3627]),.i2(intermediate_reg_0[3626]),.o(intermediate_reg_1[1813]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3625]),.i2(intermediate_reg_0[3624]),.o(intermediate_reg_1[1812])); 
mux_module mux_module_inst_1_1486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3623]),.i2(intermediate_reg_0[3622]),.o(intermediate_reg_1[1811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3621]),.i2(intermediate_reg_0[3620]),.o(intermediate_reg_1[1810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3619]),.i2(intermediate_reg_0[3618]),.o(intermediate_reg_1[1809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3617]),.i2(intermediate_reg_0[3616]),.o(intermediate_reg_1[1808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3615]),.i2(intermediate_reg_0[3614]),.o(intermediate_reg_1[1807]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3613]),.i2(intermediate_reg_0[3612]),.o(intermediate_reg_1[1806])); 
xor_module xor_module_inst_1_1492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3611]),.i2(intermediate_reg_0[3610]),.o(intermediate_reg_1[1805])); 
xor_module xor_module_inst_1_1493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3609]),.i2(intermediate_reg_0[3608]),.o(intermediate_reg_1[1804])); 
xor_module xor_module_inst_1_1494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3607]),.i2(intermediate_reg_0[3606]),.o(intermediate_reg_1[1803])); 
xor_module xor_module_inst_1_1495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3605]),.i2(intermediate_reg_0[3604]),.o(intermediate_reg_1[1802])); 
mux_module mux_module_inst_1_1496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3603]),.i2(intermediate_reg_0[3602]),.o(intermediate_reg_1[1801]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3601]),.i2(intermediate_reg_0[3600]),.o(intermediate_reg_1[1800])); 
xor_module xor_module_inst_1_1498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3599]),.i2(intermediate_reg_0[3598]),.o(intermediate_reg_1[1799])); 
xor_module xor_module_inst_1_1499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3597]),.i2(intermediate_reg_0[3596]),.o(intermediate_reg_1[1798])); 
xor_module xor_module_inst_1_1500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3595]),.i2(intermediate_reg_0[3594]),.o(intermediate_reg_1[1797])); 
xor_module xor_module_inst_1_1501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3593]),.i2(intermediate_reg_0[3592]),.o(intermediate_reg_1[1796])); 
xor_module xor_module_inst_1_1502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3591]),.i2(intermediate_reg_0[3590]),.o(intermediate_reg_1[1795])); 
mux_module mux_module_inst_1_1503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3589]),.i2(intermediate_reg_0[3588]),.o(intermediate_reg_1[1794]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3587]),.i2(intermediate_reg_0[3586]),.o(intermediate_reg_1[1793])); 
xor_module xor_module_inst_1_1505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3585]),.i2(intermediate_reg_0[3584]),.o(intermediate_reg_1[1792])); 
mux_module mux_module_inst_1_1506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3583]),.i2(intermediate_reg_0[3582]),.o(intermediate_reg_1[1791]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3581]),.i2(intermediate_reg_0[3580]),.o(intermediate_reg_1[1790]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3579]),.i2(intermediate_reg_0[3578]),.o(intermediate_reg_1[1789])); 
xor_module xor_module_inst_1_1509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3577]),.i2(intermediate_reg_0[3576]),.o(intermediate_reg_1[1788])); 
xor_module xor_module_inst_1_1510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3575]),.i2(intermediate_reg_0[3574]),.o(intermediate_reg_1[1787])); 
mux_module mux_module_inst_1_1511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3573]),.i2(intermediate_reg_0[3572]),.o(intermediate_reg_1[1786]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3571]),.i2(intermediate_reg_0[3570]),.o(intermediate_reg_1[1785]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3569]),.i2(intermediate_reg_0[3568]),.o(intermediate_reg_1[1784]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3567]),.i2(intermediate_reg_0[3566]),.o(intermediate_reg_1[1783])); 
mux_module mux_module_inst_1_1515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3565]),.i2(intermediate_reg_0[3564]),.o(intermediate_reg_1[1782]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3563]),.i2(intermediate_reg_0[3562]),.o(intermediate_reg_1[1781]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3561]),.i2(intermediate_reg_0[3560]),.o(intermediate_reg_1[1780])); 
mux_module mux_module_inst_1_1518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3559]),.i2(intermediate_reg_0[3558]),.o(intermediate_reg_1[1779]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3557]),.i2(intermediate_reg_0[3556]),.o(intermediate_reg_1[1778]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3555]),.i2(intermediate_reg_0[3554]),.o(intermediate_reg_1[1777])); 
mux_module mux_module_inst_1_1521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3553]),.i2(intermediate_reg_0[3552]),.o(intermediate_reg_1[1776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3551]),.i2(intermediate_reg_0[3550]),.o(intermediate_reg_1[1775]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3549]),.i2(intermediate_reg_0[3548]),.o(intermediate_reg_1[1774]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3547]),.i2(intermediate_reg_0[3546]),.o(intermediate_reg_1[1773]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3545]),.i2(intermediate_reg_0[3544]),.o(intermediate_reg_1[1772])); 
mux_module mux_module_inst_1_1526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3543]),.i2(intermediate_reg_0[3542]),.o(intermediate_reg_1[1771]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3541]),.i2(intermediate_reg_0[3540]),.o(intermediate_reg_1[1770])); 
mux_module mux_module_inst_1_1528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3539]),.i2(intermediate_reg_0[3538]),.o(intermediate_reg_1[1769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3537]),.i2(intermediate_reg_0[3536]),.o(intermediate_reg_1[1768]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3535]),.i2(intermediate_reg_0[3534]),.o(intermediate_reg_1[1767])); 
mux_module mux_module_inst_1_1531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3533]),.i2(intermediate_reg_0[3532]),.o(intermediate_reg_1[1766]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3531]),.i2(intermediate_reg_0[3530]),.o(intermediate_reg_1[1765])); 
mux_module mux_module_inst_1_1533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3529]),.i2(intermediate_reg_0[3528]),.o(intermediate_reg_1[1764]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3527]),.i2(intermediate_reg_0[3526]),.o(intermediate_reg_1[1763]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3525]),.i2(intermediate_reg_0[3524]),.o(intermediate_reg_1[1762])); 
xor_module xor_module_inst_1_1536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3523]),.i2(intermediate_reg_0[3522]),.o(intermediate_reg_1[1761])); 
mux_module mux_module_inst_1_1537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3521]),.i2(intermediate_reg_0[3520]),.o(intermediate_reg_1[1760]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3519]),.i2(intermediate_reg_0[3518]),.o(intermediate_reg_1[1759]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3517]),.i2(intermediate_reg_0[3516]),.o(intermediate_reg_1[1758])); 
xor_module xor_module_inst_1_1540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3515]),.i2(intermediate_reg_0[3514]),.o(intermediate_reg_1[1757])); 
xor_module xor_module_inst_1_1541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3513]),.i2(intermediate_reg_0[3512]),.o(intermediate_reg_1[1756])); 
xor_module xor_module_inst_1_1542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3511]),.i2(intermediate_reg_0[3510]),.o(intermediate_reg_1[1755])); 
mux_module mux_module_inst_1_1543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3509]),.i2(intermediate_reg_0[3508]),.o(intermediate_reg_1[1754]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3507]),.i2(intermediate_reg_0[3506]),.o(intermediate_reg_1[1753])); 
xor_module xor_module_inst_1_1545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3505]),.i2(intermediate_reg_0[3504]),.o(intermediate_reg_1[1752])); 
mux_module mux_module_inst_1_1546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3503]),.i2(intermediate_reg_0[3502]),.o(intermediate_reg_1[1751]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3501]),.i2(intermediate_reg_0[3500]),.o(intermediate_reg_1[1750])); 
xor_module xor_module_inst_1_1548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3499]),.i2(intermediate_reg_0[3498]),.o(intermediate_reg_1[1749])); 
mux_module mux_module_inst_1_1549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3497]),.i2(intermediate_reg_0[3496]),.o(intermediate_reg_1[1748]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3495]),.i2(intermediate_reg_0[3494]),.o(intermediate_reg_1[1747])); 
xor_module xor_module_inst_1_1551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3493]),.i2(intermediate_reg_0[3492]),.o(intermediate_reg_1[1746])); 
mux_module mux_module_inst_1_1552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3491]),.i2(intermediate_reg_0[3490]),.o(intermediate_reg_1[1745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3489]),.i2(intermediate_reg_0[3488]),.o(intermediate_reg_1[1744]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3487]),.i2(intermediate_reg_0[3486]),.o(intermediate_reg_1[1743])); 
xor_module xor_module_inst_1_1555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3485]),.i2(intermediate_reg_0[3484]),.o(intermediate_reg_1[1742])); 
mux_module mux_module_inst_1_1556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3483]),.i2(intermediate_reg_0[3482]),.o(intermediate_reg_1[1741]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3481]),.i2(intermediate_reg_0[3480]),.o(intermediate_reg_1[1740]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3479]),.i2(intermediate_reg_0[3478]),.o(intermediate_reg_1[1739])); 
xor_module xor_module_inst_1_1559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3477]),.i2(intermediate_reg_0[3476]),.o(intermediate_reg_1[1738])); 
mux_module mux_module_inst_1_1560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3475]),.i2(intermediate_reg_0[3474]),.o(intermediate_reg_1[1737]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3473]),.i2(intermediate_reg_0[3472]),.o(intermediate_reg_1[1736]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3471]),.i2(intermediate_reg_0[3470]),.o(intermediate_reg_1[1735]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3469]),.i2(intermediate_reg_0[3468]),.o(intermediate_reg_1[1734]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3467]),.i2(intermediate_reg_0[3466]),.o(intermediate_reg_1[1733]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3465]),.i2(intermediate_reg_0[3464]),.o(intermediate_reg_1[1732])); 
mux_module mux_module_inst_1_1566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3463]),.i2(intermediate_reg_0[3462]),.o(intermediate_reg_1[1731]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3461]),.i2(intermediate_reg_0[3460]),.o(intermediate_reg_1[1730]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3459]),.i2(intermediate_reg_0[3458]),.o(intermediate_reg_1[1729]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3457]),.i2(intermediate_reg_0[3456]),.o(intermediate_reg_1[1728])); 
xor_module xor_module_inst_1_1570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3455]),.i2(intermediate_reg_0[3454]),.o(intermediate_reg_1[1727])); 
mux_module mux_module_inst_1_1571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3453]),.i2(intermediate_reg_0[3452]),.o(intermediate_reg_1[1726]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3451]),.i2(intermediate_reg_0[3450]),.o(intermediate_reg_1[1725])); 
xor_module xor_module_inst_1_1573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3449]),.i2(intermediate_reg_0[3448]),.o(intermediate_reg_1[1724])); 
xor_module xor_module_inst_1_1574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3447]),.i2(intermediate_reg_0[3446]),.o(intermediate_reg_1[1723])); 
mux_module mux_module_inst_1_1575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3445]),.i2(intermediate_reg_0[3444]),.o(intermediate_reg_1[1722]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3443]),.i2(intermediate_reg_0[3442]),.o(intermediate_reg_1[1721]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3441]),.i2(intermediate_reg_0[3440]),.o(intermediate_reg_1[1720])); 
xor_module xor_module_inst_1_1578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3439]),.i2(intermediate_reg_0[3438]),.o(intermediate_reg_1[1719])); 
xor_module xor_module_inst_1_1579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3437]),.i2(intermediate_reg_0[3436]),.o(intermediate_reg_1[1718])); 
mux_module mux_module_inst_1_1580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3435]),.i2(intermediate_reg_0[3434]),.o(intermediate_reg_1[1717]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3433]),.i2(intermediate_reg_0[3432]),.o(intermediate_reg_1[1716]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3431]),.i2(intermediate_reg_0[3430]),.o(intermediate_reg_1[1715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3429]),.i2(intermediate_reg_0[3428]),.o(intermediate_reg_1[1714]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3427]),.i2(intermediate_reg_0[3426]),.o(intermediate_reg_1[1713])); 
xor_module xor_module_inst_1_1585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3425]),.i2(intermediate_reg_0[3424]),.o(intermediate_reg_1[1712])); 
mux_module mux_module_inst_1_1586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3423]),.i2(intermediate_reg_0[3422]),.o(intermediate_reg_1[1711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3421]),.i2(intermediate_reg_0[3420]),.o(intermediate_reg_1[1710]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3419]),.i2(intermediate_reg_0[3418]),.o(intermediate_reg_1[1709])); 
xor_module xor_module_inst_1_1589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3417]),.i2(intermediate_reg_0[3416]),.o(intermediate_reg_1[1708])); 
mux_module mux_module_inst_1_1590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3415]),.i2(intermediate_reg_0[3414]),.o(intermediate_reg_1[1707]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3413]),.i2(intermediate_reg_0[3412]),.o(intermediate_reg_1[1706])); 
mux_module mux_module_inst_1_1592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3411]),.i2(intermediate_reg_0[3410]),.o(intermediate_reg_1[1705]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3409]),.i2(intermediate_reg_0[3408]),.o(intermediate_reg_1[1704]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3407]),.i2(intermediate_reg_0[3406]),.o(intermediate_reg_1[1703])); 
mux_module mux_module_inst_1_1595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3405]),.i2(intermediate_reg_0[3404]),.o(intermediate_reg_1[1702]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3403]),.i2(intermediate_reg_0[3402]),.o(intermediate_reg_1[1701])); 
mux_module mux_module_inst_1_1597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3401]),.i2(intermediate_reg_0[3400]),.o(intermediate_reg_1[1700]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3399]),.i2(intermediate_reg_0[3398]),.o(intermediate_reg_1[1699])); 
mux_module mux_module_inst_1_1599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3397]),.i2(intermediate_reg_0[3396]),.o(intermediate_reg_1[1698]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3395]),.i2(intermediate_reg_0[3394]),.o(intermediate_reg_1[1697])); 
xor_module xor_module_inst_1_1601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3393]),.i2(intermediate_reg_0[3392]),.o(intermediate_reg_1[1696])); 
mux_module mux_module_inst_1_1602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3391]),.i2(intermediate_reg_0[3390]),.o(intermediate_reg_1[1695]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3389]),.i2(intermediate_reg_0[3388]),.o(intermediate_reg_1[1694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3387]),.i2(intermediate_reg_0[3386]),.o(intermediate_reg_1[1693]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3385]),.i2(intermediate_reg_0[3384]),.o(intermediate_reg_1[1692])); 
xor_module xor_module_inst_1_1606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3383]),.i2(intermediate_reg_0[3382]),.o(intermediate_reg_1[1691])); 
mux_module mux_module_inst_1_1607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3381]),.i2(intermediate_reg_0[3380]),.o(intermediate_reg_1[1690]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3379]),.i2(intermediate_reg_0[3378]),.o(intermediate_reg_1[1689]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3377]),.i2(intermediate_reg_0[3376]),.o(intermediate_reg_1[1688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3375]),.i2(intermediate_reg_0[3374]),.o(intermediate_reg_1[1687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3373]),.i2(intermediate_reg_0[3372]),.o(intermediate_reg_1[1686]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3371]),.i2(intermediate_reg_0[3370]),.o(intermediate_reg_1[1685])); 
mux_module mux_module_inst_1_1613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3369]),.i2(intermediate_reg_0[3368]),.o(intermediate_reg_1[1684]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3367]),.i2(intermediate_reg_0[3366]),.o(intermediate_reg_1[1683])); 
mux_module mux_module_inst_1_1615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3365]),.i2(intermediate_reg_0[3364]),.o(intermediate_reg_1[1682]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3363]),.i2(intermediate_reg_0[3362]),.o(intermediate_reg_1[1681])); 
xor_module xor_module_inst_1_1617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3361]),.i2(intermediate_reg_0[3360]),.o(intermediate_reg_1[1680])); 
xor_module xor_module_inst_1_1618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3359]),.i2(intermediate_reg_0[3358]),.o(intermediate_reg_1[1679])); 
xor_module xor_module_inst_1_1619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3357]),.i2(intermediate_reg_0[3356]),.o(intermediate_reg_1[1678])); 
xor_module xor_module_inst_1_1620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3355]),.i2(intermediate_reg_0[3354]),.o(intermediate_reg_1[1677])); 
xor_module xor_module_inst_1_1621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3353]),.i2(intermediate_reg_0[3352]),.o(intermediate_reg_1[1676])); 
xor_module xor_module_inst_1_1622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3351]),.i2(intermediate_reg_0[3350]),.o(intermediate_reg_1[1675])); 
xor_module xor_module_inst_1_1623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3349]),.i2(intermediate_reg_0[3348]),.o(intermediate_reg_1[1674])); 
mux_module mux_module_inst_1_1624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3347]),.i2(intermediate_reg_0[3346]),.o(intermediate_reg_1[1673]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3345]),.i2(intermediate_reg_0[3344]),.o(intermediate_reg_1[1672])); 
xor_module xor_module_inst_1_1626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3343]),.i2(intermediate_reg_0[3342]),.o(intermediate_reg_1[1671])); 
mux_module mux_module_inst_1_1627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3341]),.i2(intermediate_reg_0[3340]),.o(intermediate_reg_1[1670]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3339]),.i2(intermediate_reg_0[3338]),.o(intermediate_reg_1[1669]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3337]),.i2(intermediate_reg_0[3336]),.o(intermediate_reg_1[1668]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3335]),.i2(intermediate_reg_0[3334]),.o(intermediate_reg_1[1667]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3333]),.i2(intermediate_reg_0[3332]),.o(intermediate_reg_1[1666])); 
xor_module xor_module_inst_1_1632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3331]),.i2(intermediate_reg_0[3330]),.o(intermediate_reg_1[1665])); 
mux_module mux_module_inst_1_1633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3329]),.i2(intermediate_reg_0[3328]),.o(intermediate_reg_1[1664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3327]),.i2(intermediate_reg_0[3326]),.o(intermediate_reg_1[1663]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3325]),.i2(intermediate_reg_0[3324]),.o(intermediate_reg_1[1662])); 
mux_module mux_module_inst_1_1636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3323]),.i2(intermediate_reg_0[3322]),.o(intermediate_reg_1[1661]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3321]),.i2(intermediate_reg_0[3320]),.o(intermediate_reg_1[1660]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3319]),.i2(intermediate_reg_0[3318]),.o(intermediate_reg_1[1659]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3317]),.i2(intermediate_reg_0[3316]),.o(intermediate_reg_1[1658]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3315]),.i2(intermediate_reg_0[3314]),.o(intermediate_reg_1[1657])); 
mux_module mux_module_inst_1_1641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3313]),.i2(intermediate_reg_0[3312]),.o(intermediate_reg_1[1656]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3311]),.i2(intermediate_reg_0[3310]),.o(intermediate_reg_1[1655])); 
mux_module mux_module_inst_1_1643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3309]),.i2(intermediate_reg_0[3308]),.o(intermediate_reg_1[1654]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3307]),.i2(intermediate_reg_0[3306]),.o(intermediate_reg_1[1653])); 
mux_module mux_module_inst_1_1645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3305]),.i2(intermediate_reg_0[3304]),.o(intermediate_reg_1[1652]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3303]),.i2(intermediate_reg_0[3302]),.o(intermediate_reg_1[1651])); 
mux_module mux_module_inst_1_1647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3301]),.i2(intermediate_reg_0[3300]),.o(intermediate_reg_1[1650]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3299]),.i2(intermediate_reg_0[3298]),.o(intermediate_reg_1[1649])); 
mux_module mux_module_inst_1_1649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3297]),.i2(intermediate_reg_0[3296]),.o(intermediate_reg_1[1648]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3295]),.i2(intermediate_reg_0[3294]),.o(intermediate_reg_1[1647])); 
mux_module mux_module_inst_1_1651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3293]),.i2(intermediate_reg_0[3292]),.o(intermediate_reg_1[1646]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3291]),.i2(intermediate_reg_0[3290]),.o(intermediate_reg_1[1645]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3289]),.i2(intermediate_reg_0[3288]),.o(intermediate_reg_1[1644])); 
mux_module mux_module_inst_1_1654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3287]),.i2(intermediate_reg_0[3286]),.o(intermediate_reg_1[1643]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3285]),.i2(intermediate_reg_0[3284]),.o(intermediate_reg_1[1642])); 
mux_module mux_module_inst_1_1656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3283]),.i2(intermediate_reg_0[3282]),.o(intermediate_reg_1[1641]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3281]),.i2(intermediate_reg_0[3280]),.o(intermediate_reg_1[1640])); 
mux_module mux_module_inst_1_1658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3279]),.i2(intermediate_reg_0[3278]),.o(intermediate_reg_1[1639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3277]),.i2(intermediate_reg_0[3276]),.o(intermediate_reg_1[1638]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3275]),.i2(intermediate_reg_0[3274]),.o(intermediate_reg_1[1637]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3273]),.i2(intermediate_reg_0[3272]),.o(intermediate_reg_1[1636])); 
xor_module xor_module_inst_1_1662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3271]),.i2(intermediate_reg_0[3270]),.o(intermediate_reg_1[1635])); 
xor_module xor_module_inst_1_1663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3269]),.i2(intermediate_reg_0[3268]),.o(intermediate_reg_1[1634])); 
mux_module mux_module_inst_1_1664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3267]),.i2(intermediate_reg_0[3266]),.o(intermediate_reg_1[1633]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3265]),.i2(intermediate_reg_0[3264]),.o(intermediate_reg_1[1632])); 
xor_module xor_module_inst_1_1666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3263]),.i2(intermediate_reg_0[3262]),.o(intermediate_reg_1[1631])); 
xor_module xor_module_inst_1_1667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3261]),.i2(intermediate_reg_0[3260]),.o(intermediate_reg_1[1630])); 
mux_module mux_module_inst_1_1668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3259]),.i2(intermediate_reg_0[3258]),.o(intermediate_reg_1[1629]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3257]),.i2(intermediate_reg_0[3256]),.o(intermediate_reg_1[1628]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3255]),.i2(intermediate_reg_0[3254]),.o(intermediate_reg_1[1627]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3253]),.i2(intermediate_reg_0[3252]),.o(intermediate_reg_1[1626]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3251]),.i2(intermediate_reg_0[3250]),.o(intermediate_reg_1[1625])); 
xor_module xor_module_inst_1_1673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3249]),.i2(intermediate_reg_0[3248]),.o(intermediate_reg_1[1624])); 
xor_module xor_module_inst_1_1674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3247]),.i2(intermediate_reg_0[3246]),.o(intermediate_reg_1[1623])); 
xor_module xor_module_inst_1_1675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3245]),.i2(intermediate_reg_0[3244]),.o(intermediate_reg_1[1622])); 
xor_module xor_module_inst_1_1676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3243]),.i2(intermediate_reg_0[3242]),.o(intermediate_reg_1[1621])); 
mux_module mux_module_inst_1_1677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3241]),.i2(intermediate_reg_0[3240]),.o(intermediate_reg_1[1620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3239]),.i2(intermediate_reg_0[3238]),.o(intermediate_reg_1[1619]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3237]),.i2(intermediate_reg_0[3236]),.o(intermediate_reg_1[1618])); 
xor_module xor_module_inst_1_1680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3235]),.i2(intermediate_reg_0[3234]),.o(intermediate_reg_1[1617])); 
mux_module mux_module_inst_1_1681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3233]),.i2(intermediate_reg_0[3232]),.o(intermediate_reg_1[1616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3231]),.i2(intermediate_reg_0[3230]),.o(intermediate_reg_1[1615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3229]),.i2(intermediate_reg_0[3228]),.o(intermediate_reg_1[1614]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3227]),.i2(intermediate_reg_0[3226]),.o(intermediate_reg_1[1613])); 
mux_module mux_module_inst_1_1685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3225]),.i2(intermediate_reg_0[3224]),.o(intermediate_reg_1[1612]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3223]),.i2(intermediate_reg_0[3222]),.o(intermediate_reg_1[1611])); 
mux_module mux_module_inst_1_1687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3221]),.i2(intermediate_reg_0[3220]),.o(intermediate_reg_1[1610]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3219]),.i2(intermediate_reg_0[3218]),.o(intermediate_reg_1[1609])); 
mux_module mux_module_inst_1_1689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3217]),.i2(intermediate_reg_0[3216]),.o(intermediate_reg_1[1608]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3215]),.i2(intermediate_reg_0[3214]),.o(intermediate_reg_1[1607])); 
mux_module mux_module_inst_1_1691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3213]),.i2(intermediate_reg_0[3212]),.o(intermediate_reg_1[1606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3211]),.i2(intermediate_reg_0[3210]),.o(intermediate_reg_1[1605]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3209]),.i2(intermediate_reg_0[3208]),.o(intermediate_reg_1[1604])); 
mux_module mux_module_inst_1_1694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3207]),.i2(intermediate_reg_0[3206]),.o(intermediate_reg_1[1603]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3205]),.i2(intermediate_reg_0[3204]),.o(intermediate_reg_1[1602])); 
mux_module mux_module_inst_1_1696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3203]),.i2(intermediate_reg_0[3202]),.o(intermediate_reg_1[1601]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3201]),.i2(intermediate_reg_0[3200]),.o(intermediate_reg_1[1600])); 
xor_module xor_module_inst_1_1698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3199]),.i2(intermediate_reg_0[3198]),.o(intermediate_reg_1[1599])); 
xor_module xor_module_inst_1_1699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3197]),.i2(intermediate_reg_0[3196]),.o(intermediate_reg_1[1598])); 
xor_module xor_module_inst_1_1700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3195]),.i2(intermediate_reg_0[3194]),.o(intermediate_reg_1[1597])); 
xor_module xor_module_inst_1_1701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3193]),.i2(intermediate_reg_0[3192]),.o(intermediate_reg_1[1596])); 
xor_module xor_module_inst_1_1702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3191]),.i2(intermediate_reg_0[3190]),.o(intermediate_reg_1[1595])); 
mux_module mux_module_inst_1_1703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3189]),.i2(intermediate_reg_0[3188]),.o(intermediate_reg_1[1594]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3187]),.i2(intermediate_reg_0[3186]),.o(intermediate_reg_1[1593])); 
mux_module mux_module_inst_1_1705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3185]),.i2(intermediate_reg_0[3184]),.o(intermediate_reg_1[1592]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3183]),.i2(intermediate_reg_0[3182]),.o(intermediate_reg_1[1591]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3181]),.i2(intermediate_reg_0[3180]),.o(intermediate_reg_1[1590]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3179]),.i2(intermediate_reg_0[3178]),.o(intermediate_reg_1[1589]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3177]),.i2(intermediate_reg_0[3176]),.o(intermediate_reg_1[1588]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3175]),.i2(intermediate_reg_0[3174]),.o(intermediate_reg_1[1587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3173]),.i2(intermediate_reg_0[3172]),.o(intermediate_reg_1[1586]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3171]),.i2(intermediate_reg_0[3170]),.o(intermediate_reg_1[1585])); 
xor_module xor_module_inst_1_1713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3169]),.i2(intermediate_reg_0[3168]),.o(intermediate_reg_1[1584])); 
mux_module mux_module_inst_1_1714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3167]),.i2(intermediate_reg_0[3166]),.o(intermediate_reg_1[1583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3165]),.i2(intermediate_reg_0[3164]),.o(intermediate_reg_1[1582]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3163]),.i2(intermediate_reg_0[3162]),.o(intermediate_reg_1[1581])); 
xor_module xor_module_inst_1_1717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3161]),.i2(intermediate_reg_0[3160]),.o(intermediate_reg_1[1580])); 
xor_module xor_module_inst_1_1718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3159]),.i2(intermediate_reg_0[3158]),.o(intermediate_reg_1[1579])); 
mux_module mux_module_inst_1_1719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3157]),.i2(intermediate_reg_0[3156]),.o(intermediate_reg_1[1578]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3155]),.i2(intermediate_reg_0[3154]),.o(intermediate_reg_1[1577])); 
mux_module mux_module_inst_1_1721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3153]),.i2(intermediate_reg_0[3152]),.o(intermediate_reg_1[1576]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3151]),.i2(intermediate_reg_0[3150]),.o(intermediate_reg_1[1575])); 
mux_module mux_module_inst_1_1723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3149]),.i2(intermediate_reg_0[3148]),.o(intermediate_reg_1[1574]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3147]),.i2(intermediate_reg_0[3146]),.o(intermediate_reg_1[1573])); 
xor_module xor_module_inst_1_1725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3145]),.i2(intermediate_reg_0[3144]),.o(intermediate_reg_1[1572])); 
xor_module xor_module_inst_1_1726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3143]),.i2(intermediate_reg_0[3142]),.o(intermediate_reg_1[1571])); 
xor_module xor_module_inst_1_1727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3141]),.i2(intermediate_reg_0[3140]),.o(intermediate_reg_1[1570])); 
mux_module mux_module_inst_1_1728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3139]),.i2(intermediate_reg_0[3138]),.o(intermediate_reg_1[1569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3137]),.i2(intermediate_reg_0[3136]),.o(intermediate_reg_1[1568]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3135]),.i2(intermediate_reg_0[3134]),.o(intermediate_reg_1[1567])); 
xor_module xor_module_inst_1_1731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3133]),.i2(intermediate_reg_0[3132]),.o(intermediate_reg_1[1566])); 
xor_module xor_module_inst_1_1732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3131]),.i2(intermediate_reg_0[3130]),.o(intermediate_reg_1[1565])); 
mux_module mux_module_inst_1_1733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3129]),.i2(intermediate_reg_0[3128]),.o(intermediate_reg_1[1564]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3127]),.i2(intermediate_reg_0[3126]),.o(intermediate_reg_1[1563]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3125]),.i2(intermediate_reg_0[3124]),.o(intermediate_reg_1[1562]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3123]),.i2(intermediate_reg_0[3122]),.o(intermediate_reg_1[1561])); 
mux_module mux_module_inst_1_1737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3121]),.i2(intermediate_reg_0[3120]),.o(intermediate_reg_1[1560]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3119]),.i2(intermediate_reg_0[3118]),.o(intermediate_reg_1[1559]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3117]),.i2(intermediate_reg_0[3116]),.o(intermediate_reg_1[1558]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3115]),.i2(intermediate_reg_0[3114]),.o(intermediate_reg_1[1557])); 
xor_module xor_module_inst_1_1741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3113]),.i2(intermediate_reg_0[3112]),.o(intermediate_reg_1[1556])); 
xor_module xor_module_inst_1_1742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3111]),.i2(intermediate_reg_0[3110]),.o(intermediate_reg_1[1555])); 
mux_module mux_module_inst_1_1743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3109]),.i2(intermediate_reg_0[3108]),.o(intermediate_reg_1[1554]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3107]),.i2(intermediate_reg_0[3106]),.o(intermediate_reg_1[1553])); 
xor_module xor_module_inst_1_1745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3105]),.i2(intermediate_reg_0[3104]),.o(intermediate_reg_1[1552])); 
mux_module mux_module_inst_1_1746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3103]),.i2(intermediate_reg_0[3102]),.o(intermediate_reg_1[1551]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3101]),.i2(intermediate_reg_0[3100]),.o(intermediate_reg_1[1550])); 
xor_module xor_module_inst_1_1748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3099]),.i2(intermediate_reg_0[3098]),.o(intermediate_reg_1[1549])); 
xor_module xor_module_inst_1_1749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3097]),.i2(intermediate_reg_0[3096]),.o(intermediate_reg_1[1548])); 
mux_module mux_module_inst_1_1750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3095]),.i2(intermediate_reg_0[3094]),.o(intermediate_reg_1[1547]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3093]),.i2(intermediate_reg_0[3092]),.o(intermediate_reg_1[1546])); 
mux_module mux_module_inst_1_1752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3091]),.i2(intermediate_reg_0[3090]),.o(intermediate_reg_1[1545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3089]),.i2(intermediate_reg_0[3088]),.o(intermediate_reg_1[1544]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3087]),.i2(intermediate_reg_0[3086]),.o(intermediate_reg_1[1543])); 
xor_module xor_module_inst_1_1755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3085]),.i2(intermediate_reg_0[3084]),.o(intermediate_reg_1[1542])); 
mux_module mux_module_inst_1_1756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3083]),.i2(intermediate_reg_0[3082]),.o(intermediate_reg_1[1541]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3081]),.i2(intermediate_reg_0[3080]),.o(intermediate_reg_1[1540])); 
mux_module mux_module_inst_1_1758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3079]),.i2(intermediate_reg_0[3078]),.o(intermediate_reg_1[1539]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3077]),.i2(intermediate_reg_0[3076]),.o(intermediate_reg_1[1538])); 
xor_module xor_module_inst_1_1760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3075]),.i2(intermediate_reg_0[3074]),.o(intermediate_reg_1[1537])); 
xor_module xor_module_inst_1_1761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3073]),.i2(intermediate_reg_0[3072]),.o(intermediate_reg_1[1536])); 
xor_module xor_module_inst_1_1762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3071]),.i2(intermediate_reg_0[3070]),.o(intermediate_reg_1[1535])); 
xor_module xor_module_inst_1_1763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3069]),.i2(intermediate_reg_0[3068]),.o(intermediate_reg_1[1534])); 
xor_module xor_module_inst_1_1764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3067]),.i2(intermediate_reg_0[3066]),.o(intermediate_reg_1[1533])); 
xor_module xor_module_inst_1_1765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3065]),.i2(intermediate_reg_0[3064]),.o(intermediate_reg_1[1532])); 
xor_module xor_module_inst_1_1766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3063]),.i2(intermediate_reg_0[3062]),.o(intermediate_reg_1[1531])); 
mux_module mux_module_inst_1_1767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3061]),.i2(intermediate_reg_0[3060]),.o(intermediate_reg_1[1530]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3059]),.i2(intermediate_reg_0[3058]),.o(intermediate_reg_1[1529]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3057]),.i2(intermediate_reg_0[3056]),.o(intermediate_reg_1[1528])); 
xor_module xor_module_inst_1_1770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3055]),.i2(intermediate_reg_0[3054]),.o(intermediate_reg_1[1527])); 
mux_module mux_module_inst_1_1771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3053]),.i2(intermediate_reg_0[3052]),.o(intermediate_reg_1[1526]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3051]),.i2(intermediate_reg_0[3050]),.o(intermediate_reg_1[1525]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3049]),.i2(intermediate_reg_0[3048]),.o(intermediate_reg_1[1524])); 
mux_module mux_module_inst_1_1774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3047]),.i2(intermediate_reg_0[3046]),.o(intermediate_reg_1[1523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3045]),.i2(intermediate_reg_0[3044]),.o(intermediate_reg_1[1522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3043]),.i2(intermediate_reg_0[3042]),.o(intermediate_reg_1[1521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3041]),.i2(intermediate_reg_0[3040]),.o(intermediate_reg_1[1520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3039]),.i2(intermediate_reg_0[3038]),.o(intermediate_reg_1[1519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3037]),.i2(intermediate_reg_0[3036]),.o(intermediate_reg_1[1518]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3035]),.i2(intermediate_reg_0[3034]),.o(intermediate_reg_1[1517]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3033]),.i2(intermediate_reg_0[3032]),.o(intermediate_reg_1[1516]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3031]),.i2(intermediate_reg_0[3030]),.o(intermediate_reg_1[1515])); 
mux_module mux_module_inst_1_1783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3029]),.i2(intermediate_reg_0[3028]),.o(intermediate_reg_1[1514]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3027]),.i2(intermediate_reg_0[3026]),.o(intermediate_reg_1[1513]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3025]),.i2(intermediate_reg_0[3024]),.o(intermediate_reg_1[1512])); 
xor_module xor_module_inst_1_1786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3023]),.i2(intermediate_reg_0[3022]),.o(intermediate_reg_1[1511])); 
mux_module mux_module_inst_1_1787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3021]),.i2(intermediate_reg_0[3020]),.o(intermediate_reg_1[1510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3019]),.i2(intermediate_reg_0[3018]),.o(intermediate_reg_1[1509]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3017]),.i2(intermediate_reg_0[3016]),.o(intermediate_reg_1[1508])); 
mux_module mux_module_inst_1_1790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3015]),.i2(intermediate_reg_0[3014]),.o(intermediate_reg_1[1507]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3013]),.i2(intermediate_reg_0[3012]),.o(intermediate_reg_1[1506])); 
mux_module mux_module_inst_1_1792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3011]),.i2(intermediate_reg_0[3010]),.o(intermediate_reg_1[1505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3009]),.i2(intermediate_reg_0[3008]),.o(intermediate_reg_1[1504]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3007]),.i2(intermediate_reg_0[3006]),.o(intermediate_reg_1[1503])); 
xor_module xor_module_inst_1_1795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3005]),.i2(intermediate_reg_0[3004]),.o(intermediate_reg_1[1502])); 
xor_module xor_module_inst_1_1796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3003]),.i2(intermediate_reg_0[3002]),.o(intermediate_reg_1[1501])); 
mux_module mux_module_inst_1_1797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3001]),.i2(intermediate_reg_0[3000]),.o(intermediate_reg_1[1500]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2999]),.i2(intermediate_reg_0[2998]),.o(intermediate_reg_1[1499])); 
xor_module xor_module_inst_1_1799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2997]),.i2(intermediate_reg_0[2996]),.o(intermediate_reg_1[1498])); 
xor_module xor_module_inst_1_1800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2995]),.i2(intermediate_reg_0[2994]),.o(intermediate_reg_1[1497])); 
mux_module mux_module_inst_1_1801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2993]),.i2(intermediate_reg_0[2992]),.o(intermediate_reg_1[1496]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2991]),.i2(intermediate_reg_0[2990]),.o(intermediate_reg_1[1495]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2989]),.i2(intermediate_reg_0[2988]),.o(intermediate_reg_1[1494])); 
xor_module xor_module_inst_1_1804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2987]),.i2(intermediate_reg_0[2986]),.o(intermediate_reg_1[1493])); 
mux_module mux_module_inst_1_1805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2985]),.i2(intermediate_reg_0[2984]),.o(intermediate_reg_1[1492]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2983]),.i2(intermediate_reg_0[2982]),.o(intermediate_reg_1[1491])); 
mux_module mux_module_inst_1_1807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2981]),.i2(intermediate_reg_0[2980]),.o(intermediate_reg_1[1490]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2979]),.i2(intermediate_reg_0[2978]),.o(intermediate_reg_1[1489]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2977]),.i2(intermediate_reg_0[2976]),.o(intermediate_reg_1[1488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2975]),.i2(intermediate_reg_0[2974]),.o(intermediate_reg_1[1487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2973]),.i2(intermediate_reg_0[2972]),.o(intermediate_reg_1[1486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2971]),.i2(intermediate_reg_0[2970]),.o(intermediate_reg_1[1485]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2969]),.i2(intermediate_reg_0[2968]),.o(intermediate_reg_1[1484])); 
xor_module xor_module_inst_1_1814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2967]),.i2(intermediate_reg_0[2966]),.o(intermediate_reg_1[1483])); 
xor_module xor_module_inst_1_1815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2965]),.i2(intermediate_reg_0[2964]),.o(intermediate_reg_1[1482])); 
xor_module xor_module_inst_1_1816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2963]),.i2(intermediate_reg_0[2962]),.o(intermediate_reg_1[1481])); 
xor_module xor_module_inst_1_1817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2961]),.i2(intermediate_reg_0[2960]),.o(intermediate_reg_1[1480])); 
mux_module mux_module_inst_1_1818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2959]),.i2(intermediate_reg_0[2958]),.o(intermediate_reg_1[1479]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2957]),.i2(intermediate_reg_0[2956]),.o(intermediate_reg_1[1478])); 
xor_module xor_module_inst_1_1820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2955]),.i2(intermediate_reg_0[2954]),.o(intermediate_reg_1[1477])); 
xor_module xor_module_inst_1_1821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2953]),.i2(intermediate_reg_0[2952]),.o(intermediate_reg_1[1476])); 
xor_module xor_module_inst_1_1822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2951]),.i2(intermediate_reg_0[2950]),.o(intermediate_reg_1[1475])); 
xor_module xor_module_inst_1_1823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2949]),.i2(intermediate_reg_0[2948]),.o(intermediate_reg_1[1474])); 
mux_module mux_module_inst_1_1824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2947]),.i2(intermediate_reg_0[2946]),.o(intermediate_reg_1[1473]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2945]),.i2(intermediate_reg_0[2944]),.o(intermediate_reg_1[1472]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2943]),.i2(intermediate_reg_0[2942]),.o(intermediate_reg_1[1471]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2941]),.i2(intermediate_reg_0[2940]),.o(intermediate_reg_1[1470])); 
mux_module mux_module_inst_1_1828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2939]),.i2(intermediate_reg_0[2938]),.o(intermediate_reg_1[1469]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2937]),.i2(intermediate_reg_0[2936]),.o(intermediate_reg_1[1468])); 
mux_module mux_module_inst_1_1830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2935]),.i2(intermediate_reg_0[2934]),.o(intermediate_reg_1[1467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2933]),.i2(intermediate_reg_0[2932]),.o(intermediate_reg_1[1466]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2931]),.i2(intermediate_reg_0[2930]),.o(intermediate_reg_1[1465])); 
mux_module mux_module_inst_1_1833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2929]),.i2(intermediate_reg_0[2928]),.o(intermediate_reg_1[1464]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2927]),.i2(intermediate_reg_0[2926]),.o(intermediate_reg_1[1463])); 
mux_module mux_module_inst_1_1835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2925]),.i2(intermediate_reg_0[2924]),.o(intermediate_reg_1[1462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2923]),.i2(intermediate_reg_0[2922]),.o(intermediate_reg_1[1461]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2921]),.i2(intermediate_reg_0[2920]),.o(intermediate_reg_1[1460]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2919]),.i2(intermediate_reg_0[2918]),.o(intermediate_reg_1[1459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2917]),.i2(intermediate_reg_0[2916]),.o(intermediate_reg_1[1458]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2915]),.i2(intermediate_reg_0[2914]),.o(intermediate_reg_1[1457])); 
xor_module xor_module_inst_1_1841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2913]),.i2(intermediate_reg_0[2912]),.o(intermediate_reg_1[1456])); 
xor_module xor_module_inst_1_1842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2911]),.i2(intermediate_reg_0[2910]),.o(intermediate_reg_1[1455])); 
mux_module mux_module_inst_1_1843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2909]),.i2(intermediate_reg_0[2908]),.o(intermediate_reg_1[1454]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2907]),.i2(intermediate_reg_0[2906]),.o(intermediate_reg_1[1453])); 
mux_module mux_module_inst_1_1845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2905]),.i2(intermediate_reg_0[2904]),.o(intermediate_reg_1[1452]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2903]),.i2(intermediate_reg_0[2902]),.o(intermediate_reg_1[1451]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2901]),.i2(intermediate_reg_0[2900]),.o(intermediate_reg_1[1450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2899]),.i2(intermediate_reg_0[2898]),.o(intermediate_reg_1[1449]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2897]),.i2(intermediate_reg_0[2896]),.o(intermediate_reg_1[1448])); 
xor_module xor_module_inst_1_1850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2895]),.i2(intermediate_reg_0[2894]),.o(intermediate_reg_1[1447])); 
xor_module xor_module_inst_1_1851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2893]),.i2(intermediate_reg_0[2892]),.o(intermediate_reg_1[1446])); 
mux_module mux_module_inst_1_1852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2891]),.i2(intermediate_reg_0[2890]),.o(intermediate_reg_1[1445]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2889]),.i2(intermediate_reg_0[2888]),.o(intermediate_reg_1[1444]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2887]),.i2(intermediate_reg_0[2886]),.o(intermediate_reg_1[1443])); 
mux_module mux_module_inst_1_1855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2885]),.i2(intermediate_reg_0[2884]),.o(intermediate_reg_1[1442]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2883]),.i2(intermediate_reg_0[2882]),.o(intermediate_reg_1[1441])); 
xor_module xor_module_inst_1_1857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2881]),.i2(intermediate_reg_0[2880]),.o(intermediate_reg_1[1440])); 
mux_module mux_module_inst_1_1858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2879]),.i2(intermediate_reg_0[2878]),.o(intermediate_reg_1[1439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2877]),.i2(intermediate_reg_0[2876]),.o(intermediate_reg_1[1438]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2875]),.i2(intermediate_reg_0[2874]),.o(intermediate_reg_1[1437])); 
mux_module mux_module_inst_1_1861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2873]),.i2(intermediate_reg_0[2872]),.o(intermediate_reg_1[1436]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2871]),.i2(intermediate_reg_0[2870]),.o(intermediate_reg_1[1435]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2869]),.i2(intermediate_reg_0[2868]),.o(intermediate_reg_1[1434])); 
xor_module xor_module_inst_1_1864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2867]),.i2(intermediate_reg_0[2866]),.o(intermediate_reg_1[1433])); 
xor_module xor_module_inst_1_1865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2865]),.i2(intermediate_reg_0[2864]),.o(intermediate_reg_1[1432])); 
mux_module mux_module_inst_1_1866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2863]),.i2(intermediate_reg_0[2862]),.o(intermediate_reg_1[1431]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2861]),.i2(intermediate_reg_0[2860]),.o(intermediate_reg_1[1430])); 
mux_module mux_module_inst_1_1868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2859]),.i2(intermediate_reg_0[2858]),.o(intermediate_reg_1[1429]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2857]),.i2(intermediate_reg_0[2856]),.o(intermediate_reg_1[1428])); 
mux_module mux_module_inst_1_1870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2855]),.i2(intermediate_reg_0[2854]),.o(intermediate_reg_1[1427]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2853]),.i2(intermediate_reg_0[2852]),.o(intermediate_reg_1[1426]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2851]),.i2(intermediate_reg_0[2850]),.o(intermediate_reg_1[1425]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2849]),.i2(intermediate_reg_0[2848]),.o(intermediate_reg_1[1424]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2847]),.i2(intermediate_reg_0[2846]),.o(intermediate_reg_1[1423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2845]),.i2(intermediate_reg_0[2844]),.o(intermediate_reg_1[1422]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2843]),.i2(intermediate_reg_0[2842]),.o(intermediate_reg_1[1421]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2841]),.i2(intermediate_reg_0[2840]),.o(intermediate_reg_1[1420])); 
xor_module xor_module_inst_1_1878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2839]),.i2(intermediate_reg_0[2838]),.o(intermediate_reg_1[1419])); 
xor_module xor_module_inst_1_1879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2837]),.i2(intermediate_reg_0[2836]),.o(intermediate_reg_1[1418])); 
mux_module mux_module_inst_1_1880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2835]),.i2(intermediate_reg_0[2834]),.o(intermediate_reg_1[1417]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2833]),.i2(intermediate_reg_0[2832]),.o(intermediate_reg_1[1416])); 
mux_module mux_module_inst_1_1882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2831]),.i2(intermediate_reg_0[2830]),.o(intermediate_reg_1[1415]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2829]),.i2(intermediate_reg_0[2828]),.o(intermediate_reg_1[1414])); 
xor_module xor_module_inst_1_1884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2827]),.i2(intermediate_reg_0[2826]),.o(intermediate_reg_1[1413])); 
xor_module xor_module_inst_1_1885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2825]),.i2(intermediate_reg_0[2824]),.o(intermediate_reg_1[1412])); 
xor_module xor_module_inst_1_1886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2823]),.i2(intermediate_reg_0[2822]),.o(intermediate_reg_1[1411])); 
xor_module xor_module_inst_1_1887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2821]),.i2(intermediate_reg_0[2820]),.o(intermediate_reg_1[1410])); 
mux_module mux_module_inst_1_1888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2819]),.i2(intermediate_reg_0[2818]),.o(intermediate_reg_1[1409]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2817]),.i2(intermediate_reg_0[2816]),.o(intermediate_reg_1[1408])); 
mux_module mux_module_inst_1_1890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2815]),.i2(intermediate_reg_0[2814]),.o(intermediate_reg_1[1407]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2813]),.i2(intermediate_reg_0[2812]),.o(intermediate_reg_1[1406])); 
mux_module mux_module_inst_1_1892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2811]),.i2(intermediate_reg_0[2810]),.o(intermediate_reg_1[1405]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2809]),.i2(intermediate_reg_0[2808]),.o(intermediate_reg_1[1404])); 
mux_module mux_module_inst_1_1894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2807]),.i2(intermediate_reg_0[2806]),.o(intermediate_reg_1[1403]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2805]),.i2(intermediate_reg_0[2804]),.o(intermediate_reg_1[1402])); 
xor_module xor_module_inst_1_1896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2803]),.i2(intermediate_reg_0[2802]),.o(intermediate_reg_1[1401])); 
xor_module xor_module_inst_1_1897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2801]),.i2(intermediate_reg_0[2800]),.o(intermediate_reg_1[1400])); 
mux_module mux_module_inst_1_1898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2799]),.i2(intermediate_reg_0[2798]),.o(intermediate_reg_1[1399]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2797]),.i2(intermediate_reg_0[2796]),.o(intermediate_reg_1[1398])); 
xor_module xor_module_inst_1_1900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2795]),.i2(intermediate_reg_0[2794]),.o(intermediate_reg_1[1397])); 
xor_module xor_module_inst_1_1901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2793]),.i2(intermediate_reg_0[2792]),.o(intermediate_reg_1[1396])); 
mux_module mux_module_inst_1_1902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2791]),.i2(intermediate_reg_0[2790]),.o(intermediate_reg_1[1395]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2789]),.i2(intermediate_reg_0[2788]),.o(intermediate_reg_1[1394]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2787]),.i2(intermediate_reg_0[2786]),.o(intermediate_reg_1[1393])); 
mux_module mux_module_inst_1_1905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2785]),.i2(intermediate_reg_0[2784]),.o(intermediate_reg_1[1392]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2783]),.i2(intermediate_reg_0[2782]),.o(intermediate_reg_1[1391])); 
xor_module xor_module_inst_1_1907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2781]),.i2(intermediate_reg_0[2780]),.o(intermediate_reg_1[1390])); 
xor_module xor_module_inst_1_1908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2779]),.i2(intermediate_reg_0[2778]),.o(intermediate_reg_1[1389])); 
xor_module xor_module_inst_1_1909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2777]),.i2(intermediate_reg_0[2776]),.o(intermediate_reg_1[1388])); 
mux_module mux_module_inst_1_1910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2775]),.i2(intermediate_reg_0[2774]),.o(intermediate_reg_1[1387]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2773]),.i2(intermediate_reg_0[2772]),.o(intermediate_reg_1[1386])); 
mux_module mux_module_inst_1_1912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2771]),.i2(intermediate_reg_0[2770]),.o(intermediate_reg_1[1385]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2769]),.i2(intermediate_reg_0[2768]),.o(intermediate_reg_1[1384]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2767]),.i2(intermediate_reg_0[2766]),.o(intermediate_reg_1[1383]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2765]),.i2(intermediate_reg_0[2764]),.o(intermediate_reg_1[1382])); 
xor_module xor_module_inst_1_1916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2763]),.i2(intermediate_reg_0[2762]),.o(intermediate_reg_1[1381])); 
xor_module xor_module_inst_1_1917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2761]),.i2(intermediate_reg_0[2760]),.o(intermediate_reg_1[1380])); 
mux_module mux_module_inst_1_1918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2759]),.i2(intermediate_reg_0[2758]),.o(intermediate_reg_1[1379]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2757]),.i2(intermediate_reg_0[2756]),.o(intermediate_reg_1[1378])); 
mux_module mux_module_inst_1_1920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2755]),.i2(intermediate_reg_0[2754]),.o(intermediate_reg_1[1377]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2753]),.i2(intermediate_reg_0[2752]),.o(intermediate_reg_1[1376])); 
mux_module mux_module_inst_1_1922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2751]),.i2(intermediate_reg_0[2750]),.o(intermediate_reg_1[1375]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2749]),.i2(intermediate_reg_0[2748]),.o(intermediate_reg_1[1374])); 
mux_module mux_module_inst_1_1924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2747]),.i2(intermediate_reg_0[2746]),.o(intermediate_reg_1[1373]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2745]),.i2(intermediate_reg_0[2744]),.o(intermediate_reg_1[1372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2743]),.i2(intermediate_reg_0[2742]),.o(intermediate_reg_1[1371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2741]),.i2(intermediate_reg_0[2740]),.o(intermediate_reg_1[1370]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2739]),.i2(intermediate_reg_0[2738]),.o(intermediate_reg_1[1369])); 
mux_module mux_module_inst_1_1929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2737]),.i2(intermediate_reg_0[2736]),.o(intermediate_reg_1[1368]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2735]),.i2(intermediate_reg_0[2734]),.o(intermediate_reg_1[1367])); 
xor_module xor_module_inst_1_1931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2733]),.i2(intermediate_reg_0[2732]),.o(intermediate_reg_1[1366])); 
mux_module mux_module_inst_1_1932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2731]),.i2(intermediate_reg_0[2730]),.o(intermediate_reg_1[1365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2729]),.i2(intermediate_reg_0[2728]),.o(intermediate_reg_1[1364]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2727]),.i2(intermediate_reg_0[2726]),.o(intermediate_reg_1[1363])); 
mux_module mux_module_inst_1_1935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2725]),.i2(intermediate_reg_0[2724]),.o(intermediate_reg_1[1362]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2723]),.i2(intermediate_reg_0[2722]),.o(intermediate_reg_1[1361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2721]),.i2(intermediate_reg_0[2720]),.o(intermediate_reg_1[1360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2719]),.i2(intermediate_reg_0[2718]),.o(intermediate_reg_1[1359]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2717]),.i2(intermediate_reg_0[2716]),.o(intermediate_reg_1[1358])); 
mux_module mux_module_inst_1_1940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2715]),.i2(intermediate_reg_0[2714]),.o(intermediate_reg_1[1357]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2713]),.i2(intermediate_reg_0[2712]),.o(intermediate_reg_1[1356])); 
xor_module xor_module_inst_1_1942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2711]),.i2(intermediate_reg_0[2710]),.o(intermediate_reg_1[1355])); 
mux_module mux_module_inst_1_1943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2709]),.i2(intermediate_reg_0[2708]),.o(intermediate_reg_1[1354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2707]),.i2(intermediate_reg_0[2706]),.o(intermediate_reg_1[1353]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2705]),.i2(intermediate_reg_0[2704]),.o(intermediate_reg_1[1352])); 
mux_module mux_module_inst_1_1946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2703]),.i2(intermediate_reg_0[2702]),.o(intermediate_reg_1[1351]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2701]),.i2(intermediate_reg_0[2700]),.o(intermediate_reg_1[1350])); 
xor_module xor_module_inst_1_1948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2699]),.i2(intermediate_reg_0[2698]),.o(intermediate_reg_1[1349])); 
mux_module mux_module_inst_1_1949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2697]),.i2(intermediate_reg_0[2696]),.o(intermediate_reg_1[1348]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2695]),.i2(intermediate_reg_0[2694]),.o(intermediate_reg_1[1347]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2693]),.i2(intermediate_reg_0[2692]),.o(intermediate_reg_1[1346])); 
xor_module xor_module_inst_1_1952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2691]),.i2(intermediate_reg_0[2690]),.o(intermediate_reg_1[1345])); 
xor_module xor_module_inst_1_1953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2689]),.i2(intermediate_reg_0[2688]),.o(intermediate_reg_1[1344])); 
xor_module xor_module_inst_1_1954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2687]),.i2(intermediate_reg_0[2686]),.o(intermediate_reg_1[1343])); 
mux_module mux_module_inst_1_1955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2685]),.i2(intermediate_reg_0[2684]),.o(intermediate_reg_1[1342]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2683]),.i2(intermediate_reg_0[2682]),.o(intermediate_reg_1[1341])); 
xor_module xor_module_inst_1_1957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2681]),.i2(intermediate_reg_0[2680]),.o(intermediate_reg_1[1340])); 
xor_module xor_module_inst_1_1958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2679]),.i2(intermediate_reg_0[2678]),.o(intermediate_reg_1[1339])); 
xor_module xor_module_inst_1_1959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2677]),.i2(intermediate_reg_0[2676]),.o(intermediate_reg_1[1338])); 
mux_module mux_module_inst_1_1960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2675]),.i2(intermediate_reg_0[2674]),.o(intermediate_reg_1[1337]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2673]),.i2(intermediate_reg_0[2672]),.o(intermediate_reg_1[1336])); 
xor_module xor_module_inst_1_1962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2671]),.i2(intermediate_reg_0[2670]),.o(intermediate_reg_1[1335])); 
xor_module xor_module_inst_1_1963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2669]),.i2(intermediate_reg_0[2668]),.o(intermediate_reg_1[1334])); 
xor_module xor_module_inst_1_1964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2667]),.i2(intermediate_reg_0[2666]),.o(intermediate_reg_1[1333])); 
xor_module xor_module_inst_1_1965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2665]),.i2(intermediate_reg_0[2664]),.o(intermediate_reg_1[1332])); 
mux_module mux_module_inst_1_1966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2663]),.i2(intermediate_reg_0[2662]),.o(intermediate_reg_1[1331]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2661]),.i2(intermediate_reg_0[2660]),.o(intermediate_reg_1[1330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2659]),.i2(intermediate_reg_0[2658]),.o(intermediate_reg_1[1329]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2657]),.i2(intermediate_reg_0[2656]),.o(intermediate_reg_1[1328])); 
xor_module xor_module_inst_1_1970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2655]),.i2(intermediate_reg_0[2654]),.o(intermediate_reg_1[1327])); 
mux_module mux_module_inst_1_1971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2653]),.i2(intermediate_reg_0[2652]),.o(intermediate_reg_1[1326]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2651]),.i2(intermediate_reg_0[2650]),.o(intermediate_reg_1[1325])); 
mux_module mux_module_inst_1_1973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2649]),.i2(intermediate_reg_0[2648]),.o(intermediate_reg_1[1324]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2647]),.i2(intermediate_reg_0[2646]),.o(intermediate_reg_1[1323]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2645]),.i2(intermediate_reg_0[2644]),.o(intermediate_reg_1[1322])); 
xor_module xor_module_inst_1_1976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2643]),.i2(intermediate_reg_0[2642]),.o(intermediate_reg_1[1321])); 
xor_module xor_module_inst_1_1977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2641]),.i2(intermediate_reg_0[2640]),.o(intermediate_reg_1[1320])); 
xor_module xor_module_inst_1_1978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2639]),.i2(intermediate_reg_0[2638]),.o(intermediate_reg_1[1319])); 
mux_module mux_module_inst_1_1979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2637]),.i2(intermediate_reg_0[2636]),.o(intermediate_reg_1[1318]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2635]),.i2(intermediate_reg_0[2634]),.o(intermediate_reg_1[1317])); 
xor_module xor_module_inst_1_1981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2633]),.i2(intermediate_reg_0[2632]),.o(intermediate_reg_1[1316])); 
mux_module mux_module_inst_1_1982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2631]),.i2(intermediate_reg_0[2630]),.o(intermediate_reg_1[1315]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2629]),.i2(intermediate_reg_0[2628]),.o(intermediate_reg_1[1314])); 
mux_module mux_module_inst_1_1984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2627]),.i2(intermediate_reg_0[2626]),.o(intermediate_reg_1[1313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2625]),.i2(intermediate_reg_0[2624]),.o(intermediate_reg_1[1312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309])); 
mux_module mux_module_inst_1_1989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303])); 
mux_module mux_module_inst_1_1995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300])); 
xor_module xor_module_inst_1_1998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299])); 
xor_module xor_module_inst_1_1999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298])); 
mux_module mux_module_inst_1_2000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296])); 
xor_module xor_module_inst_1_2002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295])); 
xor_module xor_module_inst_1_2003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294])); 
mux_module mux_module_inst_1_2004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291])); 
mux_module mux_module_inst_1_2007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288])); 
xor_module xor_module_inst_1_2010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287])); 
mux_module mux_module_inst_1_2011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285])); 
mux_module mux_module_inst_1_2013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283])); 
xor_module xor_module_inst_1_2015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282])); 
mux_module mux_module_inst_1_2016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280])); 
mux_module mux_module_inst_1_2018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277])); 
xor_module xor_module_inst_1_2021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276])); 
mux_module mux_module_inst_1_2022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274])); 
mux_module mux_module_inst_1_2024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269])); 
xor_module xor_module_inst_1_2029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268])); 
mux_module mux_module_inst_1_2030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266])); 
xor_module xor_module_inst_1_2032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265])); 
mux_module mux_module_inst_1_2033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263])); 
mux_module mux_module_inst_1_2035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261])); 
xor_module xor_module_inst_1_2037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260])); 
mux_module mux_module_inst_1_2038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256])); 
xor_module xor_module_inst_1_2042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255])); 
mux_module mux_module_inst_1_2043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253])); 
xor_module xor_module_inst_1_2045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252])); 
mux_module mux_module_inst_1_2046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250])); 
xor_module xor_module_inst_1_2048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249])); 
xor_module xor_module_inst_1_2049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248])); 
xor_module xor_module_inst_1_2050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247])); 
xor_module xor_module_inst_1_2051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246])); 
xor_module xor_module_inst_1_2052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245])); 
mux_module mux_module_inst_1_2053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243])); 
mux_module mux_module_inst_1_2055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240])); 
xor_module xor_module_inst_1_2058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239])); 
mux_module mux_module_inst_1_2059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237])); 
xor_module xor_module_inst_1_2061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236])); 
xor_module xor_module_inst_1_2062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235])); 
mux_module mux_module_inst_1_2063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233])); 
mux_module mux_module_inst_1_2065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231])); 
mux_module mux_module_inst_1_2067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229])); 
xor_module xor_module_inst_1_2069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228])); 
xor_module xor_module_inst_1_2070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227])); 
xor_module xor_module_inst_1_2071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
xor_module xor_module_inst_1_2072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225])); 
mux_module mux_module_inst_1_2073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223])); 
mux_module mux_module_inst_1_2075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221])); 
mux_module mux_module_inst_1_2077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219])); 
xor_module xor_module_inst_1_2079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218])); 
mux_module mux_module_inst_1_2080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216])); 
xor_module xor_module_inst_1_2082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215])); 
xor_module xor_module_inst_1_2083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214])); 
mux_module mux_module_inst_1_2084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210])); 
xor_module xor_module_inst_1_2088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209])); 
xor_module xor_module_inst_1_2089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208])); 
xor_module xor_module_inst_1_2090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207])); 
mux_module mux_module_inst_1_2091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204])); 
xor_module xor_module_inst_1_2094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203])); 
mux_module mux_module_inst_1_2095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200])); 
xor_module xor_module_inst_1_2098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199])); 
xor_module xor_module_inst_1_2099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198])); 
xor_module xor_module_inst_1_2100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197])); 
mux_module mux_module_inst_1_2101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195])); 
xor_module xor_module_inst_1_2103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194])); 
mux_module mux_module_inst_1_2104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190])); 
xor_module xor_module_inst_1_2108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189])); 
mux_module mux_module_inst_1_2109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187])); 
xor_module xor_module_inst_1_2111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186])); 
xor_module xor_module_inst_1_2112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185])); 
mux_module mux_module_inst_1_2113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180])); 
mux_module mux_module_inst_1_2118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178])); 
xor_module xor_module_inst_1_2120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177])); 
mux_module mux_module_inst_1_2121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172])); 
mux_module mux_module_inst_1_2126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170])); 
mux_module mux_module_inst_1_2128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167])); 
xor_module xor_module_inst_1_2131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166])); 
mux_module mux_module_inst_1_2132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163])); 
xor_module xor_module_inst_1_2135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162])); 
mux_module mux_module_inst_1_2136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159])); 
mux_module mux_module_inst_1_2139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155])); 
mux_module mux_module_inst_1_2143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149])); 
xor_module xor_module_inst_1_2149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148])); 
mux_module mux_module_inst_1_2150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142])); 
xor_module xor_module_inst_1_2156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141])); 
xor_module xor_module_inst_1_2157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140])); 
xor_module xor_module_inst_1_2158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139])); 
xor_module xor_module_inst_1_2159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138])); 
mux_module mux_module_inst_1_2160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135])); 
mux_module mux_module_inst_1_2163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132])); 
mux_module mux_module_inst_1_2166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130])); 
mux_module mux_module_inst_1_2168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128])); 
mux_module mux_module_inst_1_2170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126])); 
xor_module xor_module_inst_1_2172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125])); 
xor_module xor_module_inst_1_2173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124])); 
xor_module xor_module_inst_1_2174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123])); 
mux_module mux_module_inst_1_2175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120])); 
xor_module xor_module_inst_1_2178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119])); 
xor_module xor_module_inst_1_2179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118])); 
mux_module mux_module_inst_1_2180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116])); 
mux_module mux_module_inst_1_2182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113])); 
xor_module xor_module_inst_1_2185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112])); 
xor_module xor_module_inst_1_2186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111])); 
mux_module mux_module_inst_1_2187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109])); 
xor_module xor_module_inst_1_2189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
mux_module mux_module_inst_1_2190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
xor_module xor_module_inst_1_2193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
xor_module xor_module_inst_1_2194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103])); 
mux_module mux_module_inst_1_2195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
mux_module mux_module_inst_1_2197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099])); 
mux_module mux_module_inst_1_2199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094])); 
mux_module mux_module_inst_1_2204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
mux_module mux_module_inst_1_2209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084])); 
xor_module xor_module_inst_1_2214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
mux_module mux_module_inst_1_2215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081])); 
mux_module mux_module_inst_1_2217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078])); 
mux_module mux_module_inst_1_2220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075])); 
mux_module mux_module_inst_1_2223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
mux_module mux_module_inst_1_2225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071])); 
mux_module mux_module_inst_1_2227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068])); 
xor_module xor_module_inst_1_2230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
xor_module xor_module_inst_1_2231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066])); 
mux_module mux_module_inst_1_2232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064])); 
xor_module xor_module_inst_1_2234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063])); 
mux_module mux_module_inst_1_2235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061])); 
xor_module xor_module_inst_1_2237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060])); 
xor_module xor_module_inst_1_2238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059])); 
mux_module mux_module_inst_1_2239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056])); 
mux_module mux_module_inst_1_2242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051])); 
mux_module mux_module_inst_1_2247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048])); 
xor_module xor_module_inst_1_2250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047])); 
mux_module mux_module_inst_1_2251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044])); 
xor_module xor_module_inst_1_2254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
mux_module mux_module_inst_1_2255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041])); 
mux_module mux_module_inst_1_2257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038])); 
xor_module xor_module_inst_1_2260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037])); 
xor_module xor_module_inst_1_2261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036])); 
xor_module xor_module_inst_1_2262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035])); 
mux_module mux_module_inst_1_2263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032])); 
xor_module xor_module_inst_1_2266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
mux_module mux_module_inst_1_2267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027])); 
mux_module mux_module_inst_1_2271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021])); 
xor_module xor_module_inst_1_2277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020])); 
mux_module mux_module_inst_1_2278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
mux_module mux_module_inst_1_2283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012])); 
xor_module xor_module_inst_1_2286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011])); 
mux_module mux_module_inst_1_2287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009])); 
xor_module xor_module_inst_1_2289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
xor_module xor_module_inst_1_2290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
xor_module xor_module_inst_1_2291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006])); 
mux_module mux_module_inst_1_2292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
mux_module mux_module_inst_1_2295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999])); 
xor_module xor_module_inst_1_2299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
xor_module xor_module_inst_1_2300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
mux_module mux_module_inst_1_2301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
xor_module xor_module_inst_1_2306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991])); 
mux_module mux_module_inst_1_2307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
mux_module mux_module_inst_1_2309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
xor_module xor_module_inst_1_2311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
xor_module xor_module_inst_1_2312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985])); 
xor_module xor_module_inst_1_2313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
mux_module mux_module_inst_1_2314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
xor_module xor_module_inst_1_2317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
mux_module mux_module_inst_1_2318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
xor_module xor_module_inst_1_2322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975])); 
mux_module mux_module_inst_1_2323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
xor_module xor_module_inst_1_2326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971])); 
xor_module xor_module_inst_1_2327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970])); 
mux_module mux_module_inst_1_2328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
mux_module mux_module_inst_1_2331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
mux_module mux_module_inst_1_2333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
xor_module xor_module_inst_1_2337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
mux_module mux_module_inst_1_2338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
mux_module mux_module_inst_1_2340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
xor_module xor_module_inst_1_2342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
mux_module mux_module_inst_1_2343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
xor_module xor_module_inst_1_2345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
xor_module xor_module_inst_1_2346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
xor_module xor_module_inst_1_2347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950])); 
xor_module xor_module_inst_1_2348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
mux_module mux_module_inst_1_2349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943])); 
xor_module xor_module_inst_1_2355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
xor_module xor_module_inst_1_2356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
mux_module mux_module_inst_1_2357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
xor_module xor_module_inst_1_2359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
mux_module mux_module_inst_1_2360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
xor_module xor_module_inst_1_2363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
xor_module xor_module_inst_1_2364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
mux_module mux_module_inst_1_2365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
xor_module xor_module_inst_1_2367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930])); 
mux_module mux_module_inst_1_2368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
xor_module xor_module_inst_1_2370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
mux_module mux_module_inst_1_2371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
xor_module xor_module_inst_1_2374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
mux_module mux_module_inst_1_2375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921])); 
xor_module xor_module_inst_1_2377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
xor_module xor_module_inst_1_2378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
mux_module mux_module_inst_1_2379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
mux_module mux_module_inst_1_2381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
mux_module mux_module_inst_1_2383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
mux_module mux_module_inst_1_2385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
mux_module mux_module_inst_1_2387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
mux_module mux_module_inst_1_2389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
mux_module mux_module_inst_1_2391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
xor_module xor_module_inst_1_2393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
xor_module xor_module_inst_1_2394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
xor_module xor_module_inst_1_2395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
xor_module xor_module_inst_1_2396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
mux_module mux_module_inst_1_2397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
xor_module xor_module_inst_1_2400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
xor_module xor_module_inst_1_2401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
xor_module xor_module_inst_1_2402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
mux_module mux_module_inst_1_2403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
xor_module xor_module_inst_1_2406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
xor_module xor_module_inst_1_2407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
mux_module mux_module_inst_1_2408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
xor_module xor_module_inst_1_2411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886])); 
mux_module mux_module_inst_1_2412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
xor_module xor_module_inst_1_2416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
xor_module xor_module_inst_1_2417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
xor_module xor_module_inst_1_2418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879])); 
mux_module mux_module_inst_1_2419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
mux_module mux_module_inst_1_2421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
xor_module xor_module_inst_1_2424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873])); 
mux_module mux_module_inst_1_2425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
xor_module xor_module_inst_1_2427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
xor_module xor_module_inst_1_2428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
xor_module xor_module_inst_1_2429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
mux_module mux_module_inst_1_2430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
mux_module mux_module_inst_1_2434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862])); 
xor_module xor_module_inst_1_2436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
mux_module mux_module_inst_1_2437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
xor_module xor_module_inst_1_2440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
mux_module mux_module_inst_1_2441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854])); 
mux_module mux_module_inst_1_2444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
xor_module xor_module_inst_1_2446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851])); 
mux_module mux_module_inst_1_2447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848])); 
xor_module xor_module_inst_1_2450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
xor_module xor_module_inst_1_2451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
mux_module mux_module_inst_1_2452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
mux_module mux_module_inst_1_2454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842])); 
xor_module xor_module_inst_1_2456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
xor_module xor_module_inst_1_2457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
xor_module xor_module_inst_1_2458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
xor_module xor_module_inst_1_2459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
mux_module mux_module_inst_1_2460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
xor_module xor_module_inst_1_2463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
mux_module mux_module_inst_1_2464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
mux_module mux_module_inst_1_2466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830])); 
mux_module mux_module_inst_1_2468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
mux_module mux_module_inst_1_2470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
mux_module mux_module_inst_1_2472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824])); 
mux_module mux_module_inst_1_2474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
xor_module xor_module_inst_1_2477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820])); 
mux_module mux_module_inst_1_2478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
mux_module mux_module_inst_1_2480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
xor_module xor_module_inst_1_2483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
xor_module xor_module_inst_1_2484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
mux_module mux_module_inst_1_2485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810])); 
xor_module xor_module_inst_1_2488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
mux_module mux_module_inst_1_2489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
mux_module mux_module_inst_1_2492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
xor_module xor_module_inst_1_2494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803])); 
mux_module mux_module_inst_1_2495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
xor_module xor_module_inst_1_2497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
xor_module xor_module_inst_1_2498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
mux_module mux_module_inst_1_2499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
xor_module xor_module_inst_1_2501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
xor_module xor_module_inst_1_2502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
mux_module mux_module_inst_1_2503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
mux_module mux_module_inst_1_2505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
xor_module xor_module_inst_1_2512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
mux_module mux_module_inst_1_2513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
mux_module mux_module_inst_1_2515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
xor_module xor_module_inst_1_2517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
xor_module xor_module_inst_1_2518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
xor_module xor_module_inst_1_2519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
xor_module xor_module_inst_1_2520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
mux_module mux_module_inst_1_2521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
xor_module xor_module_inst_1_2523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
xor_module xor_module_inst_1_2524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773])); 
mux_module mux_module_inst_1_2525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
mux_module mux_module_inst_1_2527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
mux_module mux_module_inst_1_2529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
xor_module xor_module_inst_1_2531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
xor_module xor_module_inst_1_2532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
xor_module xor_module_inst_1_2533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
mux_module mux_module_inst_1_2534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
mux_module mux_module_inst_1_2538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
xor_module xor_module_inst_1_2540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
mux_module mux_module_inst_1_2541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
mux_module mux_module_inst_1_2551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
xor_module xor_module_inst_1_2556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
xor_module xor_module_inst_1_2557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
xor_module xor_module_inst_1_2558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
xor_module xor_module_inst_1_2559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738])); 
mux_module mux_module_inst_1_2560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
xor_module xor_module_inst_1_2562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
mux_module mux_module_inst_1_2563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
xor_module xor_module_inst_1_2565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
mux_module mux_module_inst_1_2566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
mux_module mux_module_inst_1_2568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
mux_module mux_module_inst_1_2570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
xor_module xor_module_inst_1_2574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
xor_module xor_module_inst_1_2575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
xor_module xor_module_inst_1_2576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
xor_module xor_module_inst_1_2577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
mux_module mux_module_inst_1_2578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
xor_module xor_module_inst_1_2580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
xor_module xor_module_inst_1_2581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
mux_module mux_module_inst_1_2582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
xor_module xor_module_inst_1_2585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
mux_module mux_module_inst_1_2586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
mux_module mux_module_inst_1_2589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
xor_module xor_module_inst_1_2591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
xor_module xor_module_inst_1_2592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
xor_module xor_module_inst_1_2593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
xor_module xor_module_inst_1_2594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
xor_module xor_module_inst_1_2595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
xor_module xor_module_inst_1_2596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701])); 
xor_module xor_module_inst_1_2597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
xor_module xor_module_inst_1_2598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
xor_module xor_module_inst_1_2599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
mux_module mux_module_inst_1_2600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
mux_module mux_module_inst_1_2603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
mux_module mux_module_inst_1_2605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
mux_module mux_module_inst_1_2607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
mux_module mux_module_inst_1_2609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
xor_module xor_module_inst_1_2613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
xor_module xor_module_inst_1_2614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
mux_module mux_module_inst_1_2615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
xor_module xor_module_inst_1_2617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
mux_module mux_module_inst_1_2618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
xor_module xor_module_inst_1_2622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
mux_module mux_module_inst_1_2623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
xor_module xor_module_inst_1_2625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
xor_module xor_module_inst_1_2626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_2627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
xor_module xor_module_inst_1_2628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
xor_module xor_module_inst_1_2629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
mux_module mux_module_inst_1_2630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
xor_module xor_module_inst_1_2632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
mux_module mux_module_inst_1_2633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
mux_module mux_module_inst_1_2636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
xor_module xor_module_inst_1_2640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
mux_module mux_module_inst_1_2641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
xor_module xor_module_inst_1_2644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
xor_module xor_module_inst_1_2645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
mux_module mux_module_inst_1_2646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
xor_module xor_module_inst_1_2651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
mux_module mux_module_inst_1_2652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
mux_module mux_module_inst_1_2662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
mux_module mux_module_inst_1_2666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
mux_module mux_module_inst_1_2671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
mux_module mux_module_inst_1_2675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
mux_module mux_module_inst_1_2677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
xor_module xor_module_inst_1_2680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
xor_module xor_module_inst_1_2681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
mux_module mux_module_inst_1_2682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
mux_module mux_module_inst_1_2687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
mux_module mux_module_inst_1_2693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
xor_module xor_module_inst_1_2696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
xor_module xor_module_inst_1_2697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
mux_module mux_module_inst_1_2698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
mux_module mux_module_inst_1_2703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
xor_module xor_module_inst_1_2706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
mux_module mux_module_inst_1_2707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
xor_module xor_module_inst_1_2710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
xor_module xor_module_inst_1_2711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
xor_module xor_module_inst_1_2712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
xor_module xor_module_inst_1_2713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
xor_module xor_module_inst_1_2714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
xor_module xor_module_inst_1_2715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
mux_module mux_module_inst_1_2716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
xor_module xor_module_inst_1_2719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
xor_module xor_module_inst_1_2720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
mux_module mux_module_inst_1_2721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
mux_module mux_module_inst_1_2723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
mux_module mux_module_inst_1_2725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
xor_module xor_module_inst_1_2728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
xor_module xor_module_inst_1_2729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
xor_module xor_module_inst_1_2730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
xor_module xor_module_inst_1_2731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
xor_module xor_module_inst_1_2732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
mux_module mux_module_inst_1_2733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
mux_module mux_module_inst_1_2735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
mux_module mux_module_inst_1_2738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
xor_module xor_module_inst_1_2741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
xor_module xor_module_inst_1_2742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
xor_module xor_module_inst_1_2743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
mux_module mux_module_inst_1_2744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
mux_module mux_module_inst_1_2747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
xor_module xor_module_inst_1_2749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
xor_module xor_module_inst_1_2750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
xor_module xor_module_inst_1_2751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
xor_module xor_module_inst_1_2752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
xor_module xor_module_inst_1_2753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
mux_module mux_module_inst_1_2754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
xor_module xor_module_inst_1_2756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
xor_module xor_module_inst_1_2757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
xor_module xor_module_inst_1_2758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
xor_module xor_module_inst_1_2759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
xor_module xor_module_inst_1_2760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
xor_module xor_module_inst_1_2761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
xor_module xor_module_inst_1_2762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
mux_module mux_module_inst_1_2763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
xor_module xor_module_inst_1_2766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
xor_module xor_module_inst_1_2767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
xor_module xor_module_inst_1_2768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
mux_module mux_module_inst_1_2769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
xor_module xor_module_inst_1_2772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
xor_module xor_module_inst_1_2773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
xor_module xor_module_inst_1_2774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
xor_module xor_module_inst_1_2775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
mux_module mux_module_inst_1_2776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
xor_module xor_module_inst_1_2779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
xor_module xor_module_inst_1_2780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
mux_module mux_module_inst_1_2781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
xor_module xor_module_inst_1_2783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
xor_module xor_module_inst_1_2784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
xor_module xor_module_inst_1_2785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
xor_module xor_module_inst_1_2786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
xor_module xor_module_inst_1_2787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
xor_module xor_module_inst_1_2788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
mux_module mux_module_inst_1_2789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
xor_module xor_module_inst_1_2791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
xor_module xor_module_inst_1_2792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
xor_module xor_module_inst_1_2793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
xor_module xor_module_inst_1_2794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
mux_module mux_module_inst_1_2795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
xor_module xor_module_inst_1_2798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
mux_module mux_module_inst_1_2799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
xor_module xor_module_inst_1_2802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
mux_module mux_module_inst_1_2803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
xor_module xor_module_inst_1_2805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
mux_module mux_module_inst_1_2806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
xor_module xor_module_inst_1_2810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
xor_module xor_module_inst_1_2811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
mux_module mux_module_inst_1_2812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
xor_module xor_module_inst_1_2814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
xor_module xor_module_inst_1_2815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_2816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
xor_module xor_module_inst_1_2819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
mux_module mux_module_inst_1_2820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
xor_module xor_module_inst_1_2822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
xor_module xor_module_inst_1_2823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
mux_module mux_module_inst_1_2824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
xor_module xor_module_inst_1_2826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
mux_module mux_module_inst_1_2827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
xor_module xor_module_inst_1_2829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
xor_module xor_module_inst_1_2830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
xor_module xor_module_inst_1_2831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
xor_module xor_module_inst_1_2832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
xor_module xor_module_inst_1_2833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
mux_module mux_module_inst_1_2834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
mux_module mux_module_inst_1_2838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
mux_module mux_module_inst_1_2840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
mux_module mux_module_inst_1_2842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
xor_module xor_module_inst_1_2844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
xor_module xor_module_inst_1_2845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
mux_module mux_module_inst_1_2846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
xor_module xor_module_inst_1_2848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
mux_module mux_module_inst_1_2849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
mux_module mux_module_inst_1_2851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
mux_module mux_module_inst_1_2853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
mux_module mux_module_inst_1_2855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
xor_module xor_module_inst_1_2858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
mux_module mux_module_inst_1_2859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
mux_module mux_module_inst_1_2861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
xor_module xor_module_inst_1_2864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
mux_module mux_module_inst_1_2865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
mux_module mux_module_inst_1_2867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
mux_module mux_module_inst_1_2869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
mux_module mux_module_inst_1_2873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
mux_module mux_module_inst_1_2875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
xor_module xor_module_inst_1_2878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
mux_module mux_module_inst_1_2879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
xor_module xor_module_inst_1_2881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
xor_module xor_module_inst_1_2882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
xor_module xor_module_inst_1_2883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
xor_module xor_module_inst_1_2884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
mux_module mux_module_inst_1_2885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
xor_module xor_module_inst_1_2887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
mux_module mux_module_inst_1_2888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
mux_module mux_module_inst_1_2890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
xor_module xor_module_inst_1_2893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
mux_module mux_module_inst_1_2894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
xor_module xor_module_inst_1_2898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
xor_module xor_module_inst_1_2899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
xor_module xor_module_inst_1_2900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
mux_module mux_module_inst_1_2901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
mux_module mux_module_inst_1_2903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
mux_module mux_module_inst_1_2905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_2908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
mux_module mux_module_inst_1_2909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
mux_module mux_module_inst_1_2911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
xor_module xor_module_inst_1_2915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
xor_module xor_module_inst_1_2916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
xor_module xor_module_inst_1_2917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
xor_module xor_module_inst_1_2918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
xor_module xor_module_inst_1_2919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
xor_module xor_module_inst_1_2920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
xor_module xor_module_inst_1_2921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_2922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
mux_module mux_module_inst_1_2925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
xor_module xor_module_inst_1_2929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
mux_module mux_module_inst_1_2930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
xor_module xor_module_inst_1_2933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
mux_module mux_module_inst_1_2934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
xor_module xor_module_inst_1_2936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
mux_module mux_module_inst_1_2937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
mux_module mux_module_inst_1_2940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
xor_module xor_module_inst_1_2943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
mux_module mux_module_inst_1_2944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
xor_module xor_module_inst_1_2947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
xor_module xor_module_inst_1_2948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
xor_module xor_module_inst_1_2949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
mux_module mux_module_inst_1_2950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
mux_module mux_module_inst_1_2958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
mux_module mux_module_inst_1_2961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
mux_module mux_module_inst_1_2963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
xor_module xor_module_inst_1_2966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_2967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
xor_module xor_module_inst_1_2969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
mux_module mux_module_inst_1_2970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_2972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
mux_module mux_module_inst_1_2973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
xor_module xor_module_inst_1_2976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
xor_module xor_module_inst_1_2977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
xor_module xor_module_inst_1_2978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
mux_module mux_module_inst_1_2979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
xor_module xor_module_inst_1_2981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
mux_module mux_module_inst_1_2982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
xor_module xor_module_inst_1_2984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
xor_module xor_module_inst_1_2985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
xor_module xor_module_inst_1_2986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
xor_module xor_module_inst_1_2987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
xor_module xor_module_inst_1_2988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
mux_module mux_module_inst_1_2989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
mux_module mux_module_inst_1_2991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
xor_module xor_module_inst_1_2997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
xor_module xor_module_inst_1_2998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
mux_module mux_module_inst_1_2999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
xor_module xor_module_inst_1_3001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
mux_module mux_module_inst_1_3002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_3004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
xor_module xor_module_inst_1_3005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
xor_module xor_module_inst_1_3006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
mux_module mux_module_inst_1_3007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_3009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
xor_module xor_module_inst_1_3010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
mux_module mux_module_inst_1_3011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
xor_module xor_module_inst_1_3014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
mux_module mux_module_inst_1_3015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
mux_module mux_module_inst_1_3022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
mux_module mux_module_inst_1_3029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
xor_module xor_module_inst_1_3033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
mux_module mux_module_inst_1_3034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
mux_module mux_module_inst_1_3036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
mux_module mux_module_inst_1_3038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
mux_module mux_module_inst_1_3040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
mux_module mux_module_inst_1_3043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
xor_module xor_module_inst_1_3046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
mux_module mux_module_inst_1_3047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
mux_module mux_module_inst_1_3049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
xor_module xor_module_inst_1_3052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
xor_module xor_module_inst_1_3053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
xor_module xor_module_inst_1_3054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
xor_module xor_module_inst_1_3055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
xor_module xor_module_inst_1_3056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
mux_module mux_module_inst_1_3057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
xor_module xor_module_inst_1_3063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
xor_module xor_module_inst_1_3064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
xor_module xor_module_inst_1_3065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
mux_module mux_module_inst_1_3066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
mux_module mux_module_inst_1_3069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
xor_module xor_module_inst_1_3074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
mux_module mux_module_inst_1_3075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
mux_module mux_module_inst_1_3077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
xor_module xor_module_inst_1_3079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
xor_module xor_module_inst_1_3080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
xor_module xor_module_inst_1_3081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
mux_module mux_module_inst_1_3082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
xor_module xor_module_inst_1_3084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
mux_module mux_module_inst_1_3085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
xor_module xor_module_inst_1_3088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
xor_module xor_module_inst_1_3089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
mux_module mux_module_inst_1_3090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
mux_module mux_module_inst_1_3092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
mux_module mux_module_inst_1_3094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
mux_module mux_module_inst_1_3096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
xor_module xor_module_inst_1_3098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
xor_module xor_module_inst_1_3099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_3100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
xor_module xor_module_inst_1_3103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
mux_module mux_module_inst_1_3104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
xor_module xor_module_inst_1_3113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
mux_module mux_module_inst_1_3114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
mux_module mux_module_inst_1_3117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
mux_module mux_module_inst_1_3119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
mux_module mux_module_inst_1_3121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
xor_module xor_module_inst_1_3123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
mux_module mux_module_inst_1_3124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
xor_module xor_module_inst_1_3126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
xor_module xor_module_inst_1_3127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
xor_module xor_module_inst_1_3128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
xor_module xor_module_inst_1_3129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
mux_module mux_module_inst_1_3130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
mux_module mux_module_inst_1_3132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
xor_module xor_module_inst_1_3134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
xor_module xor_module_inst_1_3135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
xor_module xor_module_inst_1_3136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
xor_module xor_module_inst_1_3137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
mux_module mux_module_inst_1_3138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
xor_module xor_module_inst_1_3140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
mux_module mux_module_inst_1_3141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
mux_module mux_module_inst_1_3144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
xor_module xor_module_inst_1_3146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
mux_module mux_module_inst_1_3147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
xor_module xor_module_inst_1_3154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
mux_module mux_module_inst_1_3155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
mux_module mux_module_inst_1_3158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
xor_module xor_module_inst_1_3162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
xor_module xor_module_inst_1_3163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
xor_module xor_module_inst_1_3164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
mux_module mux_module_inst_1_3165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
xor_module xor_module_inst_1_3167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
mux_module mux_module_inst_1_3168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
mux_module mux_module_inst_1_3170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
mux_module mux_module_inst_1_3174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
mux_module mux_module_inst_1_3176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
mux_module mux_module_inst_1_3179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
xor_module xor_module_inst_1_3182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
mux_module mux_module_inst_1_3183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
mux_module mux_module_inst_1_3187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
xor_module xor_module_inst_1_3189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
xor_module xor_module_inst_1_3190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
mux_module mux_module_inst_1_3191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
xor_module xor_module_inst_1_3193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
mux_module mux_module_inst_1_3194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
xor_module xor_module_inst_1_3199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
xor_module xor_module_inst_1_3200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
mux_module mux_module_inst_1_3201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
xor_module xor_module_inst_1_3205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
xor_module xor_module_inst_1_3206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
mux_module mux_module_inst_1_3207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
mux_module mux_module_inst_1_3210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
mux_module mux_module_inst_1_3214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
mux_module mux_module_inst_1_3219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
mux_module mux_module_inst_1_3222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
xor_module xor_module_inst_1_3227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
mux_module mux_module_inst_1_3228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
xor_module xor_module_inst_1_3231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
xor_module xor_module_inst_1_3232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
xor_module xor_module_inst_1_3233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_3234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
mux_module mux_module_inst_1_3235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
mux_module mux_module_inst_1_3238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
xor_module xor_module_inst_1_3242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
xor_module xor_module_inst_1_3243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
xor_module xor_module_inst_1_3244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
mux_module mux_module_inst_1_3245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
mux_module mux_module_inst_1_3247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
xor_module xor_module_inst_1_3250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
mux_module mux_module_inst_1_3251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
mux_module mux_module_inst_1_3254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
mux_module mux_module_inst_1_3260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
mux_module mux_module_inst_1_3262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_3264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
mux_module mux_module_inst_1_3265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
mux_module mux_module_inst_1_3267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
mux_module mux_module_inst_1_3269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
xor_module xor_module_inst_1_3271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
xor_module xor_module_inst_1_3272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
xor_module xor_module_inst_1_3273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
mux_module mux_module_inst_1_3274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
xor_module xor_module_inst_1_3279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
xor_module xor_module_inst_1_3280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
xor_module xor_module_inst_1_3281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
mux_module mux_module_inst_1_3282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
xor_module xor_module_inst_1_3284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
xor_module xor_module_inst_1_3285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
mux_module mux_module_inst_1_3286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
mux_module mux_module_inst_1_3288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
mux_module mux_module_inst_1_3290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
xor_module xor_module_inst_1_3292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
xor_module xor_module_inst_1_3293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_3294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
mux_module mux_module_inst_1_3295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
xor_module xor_module_inst_1_3297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [3297:0] <= intermediate_reg_1; 
outp[5119:3298] <= intermediate_reg_1[1821:0] ; 
end 
endmodule 
 

module interface_12(input [6595:0] inp, output reg [835:0] outp, input clk, input reset);
reg [6595:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
wire [3297:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6595]),.i2(intermediate_reg_0[6594]),.o(intermediate_reg_1[3297]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6593]),.i2(intermediate_reg_0[6592]),.o(intermediate_reg_1[3296])); 
xor_module xor_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6591]),.i2(intermediate_reg_0[6590]),.o(intermediate_reg_1[3295])); 
xor_module xor_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6589]),.i2(intermediate_reg_0[6588]),.o(intermediate_reg_1[3294])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6587]),.i2(intermediate_reg_0[6586]),.o(intermediate_reg_1[3293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6585]),.i2(intermediate_reg_0[6584]),.o(intermediate_reg_1[3292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6583]),.i2(intermediate_reg_0[6582]),.o(intermediate_reg_1[3291]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6581]),.i2(intermediate_reg_0[6580]),.o(intermediate_reg_1[3290])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6579]),.i2(intermediate_reg_0[6578]),.o(intermediate_reg_1[3289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6577]),.i2(intermediate_reg_0[6576]),.o(intermediate_reg_1[3288]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6575]),.i2(intermediate_reg_0[6574]),.o(intermediate_reg_1[3287]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6573]),.i2(intermediate_reg_0[6572]),.o(intermediate_reg_1[3286]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6571]),.i2(intermediate_reg_0[6570]),.o(intermediate_reg_1[3285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6569]),.i2(intermediate_reg_0[6568]),.o(intermediate_reg_1[3284]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6567]),.i2(intermediate_reg_0[6566]),.o(intermediate_reg_1[3283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6565]),.i2(intermediate_reg_0[6564]),.o(intermediate_reg_1[3282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6563]),.i2(intermediate_reg_0[6562]),.o(intermediate_reg_1[3281]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6561]),.i2(intermediate_reg_0[6560]),.o(intermediate_reg_1[3280])); 
xor_module xor_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6559]),.i2(intermediate_reg_0[6558]),.o(intermediate_reg_1[3279])); 
xor_module xor_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6557]),.i2(intermediate_reg_0[6556]),.o(intermediate_reg_1[3278])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6555]),.i2(intermediate_reg_0[6554]),.o(intermediate_reg_1[3277])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6553]),.i2(intermediate_reg_0[6552]),.o(intermediate_reg_1[3276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6551]),.i2(intermediate_reg_0[6550]),.o(intermediate_reg_1[3275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6549]),.i2(intermediate_reg_0[6548]),.o(intermediate_reg_1[3274]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6547]),.i2(intermediate_reg_0[6546]),.o(intermediate_reg_1[3273]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6545]),.i2(intermediate_reg_0[6544]),.o(intermediate_reg_1[3272])); 
mux_module mux_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6543]),.i2(intermediate_reg_0[6542]),.o(intermediate_reg_1[3271]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6541]),.i2(intermediate_reg_0[6540]),.o(intermediate_reg_1[3270])); 
xor_module xor_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6539]),.i2(intermediate_reg_0[6538]),.o(intermediate_reg_1[3269])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6537]),.i2(intermediate_reg_0[6536]),.o(intermediate_reg_1[3268]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6535]),.i2(intermediate_reg_0[6534]),.o(intermediate_reg_1[3267])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6533]),.i2(intermediate_reg_0[6532]),.o(intermediate_reg_1[3266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6531]),.i2(intermediate_reg_0[6530]),.o(intermediate_reg_1[3265]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6529]),.i2(intermediate_reg_0[6528]),.o(intermediate_reg_1[3264])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6527]),.i2(intermediate_reg_0[6526]),.o(intermediate_reg_1[3263])); 
mux_module mux_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6525]),.i2(intermediate_reg_0[6524]),.o(intermediate_reg_1[3262]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6523]),.i2(intermediate_reg_0[6522]),.o(intermediate_reg_1[3261])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6521]),.i2(intermediate_reg_0[6520]),.o(intermediate_reg_1[3260])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6519]),.i2(intermediate_reg_0[6518]),.o(intermediate_reg_1[3259]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6517]),.i2(intermediate_reg_0[6516]),.o(intermediate_reg_1[3258])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6515]),.i2(intermediate_reg_0[6514]),.o(intermediate_reg_1[3257])); 
mux_module mux_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6513]),.i2(intermediate_reg_0[6512]),.o(intermediate_reg_1[3256]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6511]),.i2(intermediate_reg_0[6510]),.o(intermediate_reg_1[3255])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6509]),.i2(intermediate_reg_0[6508]),.o(intermediate_reg_1[3254])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6507]),.i2(intermediate_reg_0[6506]),.o(intermediate_reg_1[3253])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6505]),.i2(intermediate_reg_0[6504]),.o(intermediate_reg_1[3252]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6503]),.i2(intermediate_reg_0[6502]),.o(intermediate_reg_1[3251])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6501]),.i2(intermediate_reg_0[6500]),.o(intermediate_reg_1[3250])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6499]),.i2(intermediate_reg_0[6498]),.o(intermediate_reg_1[3249])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6497]),.i2(intermediate_reg_0[6496]),.o(intermediate_reg_1[3248]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6495]),.i2(intermediate_reg_0[6494]),.o(intermediate_reg_1[3247])); 
xor_module xor_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6493]),.i2(intermediate_reg_0[6492]),.o(intermediate_reg_1[3246])); 
xor_module xor_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6491]),.i2(intermediate_reg_0[6490]),.o(intermediate_reg_1[3245])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6489]),.i2(intermediate_reg_0[6488]),.o(intermediate_reg_1[3244]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6487]),.i2(intermediate_reg_0[6486]),.o(intermediate_reg_1[3243]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6485]),.i2(intermediate_reg_0[6484]),.o(intermediate_reg_1[3242])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6483]),.i2(intermediate_reg_0[6482]),.o(intermediate_reg_1[3241])); 
xor_module xor_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6481]),.i2(intermediate_reg_0[6480]),.o(intermediate_reg_1[3240])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6479]),.i2(intermediate_reg_0[6478]),.o(intermediate_reg_1[3239])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6477]),.i2(intermediate_reg_0[6476]),.o(intermediate_reg_1[3238]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6475]),.i2(intermediate_reg_0[6474]),.o(intermediate_reg_1[3237])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6473]),.i2(intermediate_reg_0[6472]),.o(intermediate_reg_1[3236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6471]),.i2(intermediate_reg_0[6470]),.o(intermediate_reg_1[3235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6469]),.i2(intermediate_reg_0[6468]),.o(intermediate_reg_1[3234]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6467]),.i2(intermediate_reg_0[6466]),.o(intermediate_reg_1[3233])); 
mux_module mux_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6465]),.i2(intermediate_reg_0[6464]),.o(intermediate_reg_1[3232]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6463]),.i2(intermediate_reg_0[6462]),.o(intermediate_reg_1[3231]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6461]),.i2(intermediate_reg_0[6460]),.o(intermediate_reg_1[3230]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6459]),.i2(intermediate_reg_0[6458]),.o(intermediate_reg_1[3229]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6457]),.i2(intermediate_reg_0[6456]),.o(intermediate_reg_1[3228])); 
xor_module xor_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6455]),.i2(intermediate_reg_0[6454]),.o(intermediate_reg_1[3227])); 
xor_module xor_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6453]),.i2(intermediate_reg_0[6452]),.o(intermediate_reg_1[3226])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6451]),.i2(intermediate_reg_0[6450]),.o(intermediate_reg_1[3225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6449]),.i2(intermediate_reg_0[6448]),.o(intermediate_reg_1[3224])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6447]),.i2(intermediate_reg_0[6446]),.o(intermediate_reg_1[3223]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6445]),.i2(intermediate_reg_0[6444]),.o(intermediate_reg_1[3222]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6443]),.i2(intermediate_reg_0[6442]),.o(intermediate_reg_1[3221])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6441]),.i2(intermediate_reg_0[6440]),.o(intermediate_reg_1[3220]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6439]),.i2(intermediate_reg_0[6438]),.o(intermediate_reg_1[3219])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6437]),.i2(intermediate_reg_0[6436]),.o(intermediate_reg_1[3218]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6435]),.i2(intermediate_reg_0[6434]),.o(intermediate_reg_1[3217])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6433]),.i2(intermediate_reg_0[6432]),.o(intermediate_reg_1[3216])); 
xor_module xor_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6431]),.i2(intermediate_reg_0[6430]),.o(intermediate_reg_1[3215])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6429]),.i2(intermediate_reg_0[6428]),.o(intermediate_reg_1[3214])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6427]),.i2(intermediate_reg_0[6426]),.o(intermediate_reg_1[3213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6425]),.i2(intermediate_reg_0[6424]),.o(intermediate_reg_1[3212]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6423]),.i2(intermediate_reg_0[6422]),.o(intermediate_reg_1[3211])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6421]),.i2(intermediate_reg_0[6420]),.o(intermediate_reg_1[3210])); 
mux_module mux_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6419]),.i2(intermediate_reg_0[6418]),.o(intermediate_reg_1[3209]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6417]),.i2(intermediate_reg_0[6416]),.o(intermediate_reg_1[3208])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6415]),.i2(intermediate_reg_0[6414]),.o(intermediate_reg_1[3207]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6413]),.i2(intermediate_reg_0[6412]),.o(intermediate_reg_1[3206])); 
xor_module xor_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6411]),.i2(intermediate_reg_0[6410]),.o(intermediate_reg_1[3205])); 
mux_module mux_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6409]),.i2(intermediate_reg_0[6408]),.o(intermediate_reg_1[3204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6407]),.i2(intermediate_reg_0[6406]),.o(intermediate_reg_1[3203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6405]),.i2(intermediate_reg_0[6404]),.o(intermediate_reg_1[3202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6403]),.i2(intermediate_reg_0[6402]),.o(intermediate_reg_1[3201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6401]),.i2(intermediate_reg_0[6400]),.o(intermediate_reg_1[3200]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6399]),.i2(intermediate_reg_0[6398]),.o(intermediate_reg_1[3199])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6397]),.i2(intermediate_reg_0[6396]),.o(intermediate_reg_1[3198])); 
mux_module mux_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6395]),.i2(intermediate_reg_0[6394]),.o(intermediate_reg_1[3197]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6393]),.i2(intermediate_reg_0[6392]),.o(intermediate_reg_1[3196])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6391]),.i2(intermediate_reg_0[6390]),.o(intermediate_reg_1[3195]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6389]),.i2(intermediate_reg_0[6388]),.o(intermediate_reg_1[3194])); 
xor_module xor_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6387]),.i2(intermediate_reg_0[6386]),.o(intermediate_reg_1[3193])); 
mux_module mux_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6385]),.i2(intermediate_reg_0[6384]),.o(intermediate_reg_1[3192]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6383]),.i2(intermediate_reg_0[6382]),.o(intermediate_reg_1[3191])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6381]),.i2(intermediate_reg_0[6380]),.o(intermediate_reg_1[3190]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6379]),.i2(intermediate_reg_0[6378]),.o(intermediate_reg_1[3189])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6377]),.i2(intermediate_reg_0[6376]),.o(intermediate_reg_1[3188])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6375]),.i2(intermediate_reg_0[6374]),.o(intermediate_reg_1[3187]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6373]),.i2(intermediate_reg_0[6372]),.o(intermediate_reg_1[3186])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6371]),.i2(intermediate_reg_0[6370]),.o(intermediate_reg_1[3185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6369]),.i2(intermediate_reg_0[6368]),.o(intermediate_reg_1[3184]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6367]),.i2(intermediate_reg_0[6366]),.o(intermediate_reg_1[3183]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6365]),.i2(intermediate_reg_0[6364]),.o(intermediate_reg_1[3182])); 
xor_module xor_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6363]),.i2(intermediate_reg_0[6362]),.o(intermediate_reg_1[3181])); 
mux_module mux_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6361]),.i2(intermediate_reg_0[6360]),.o(intermediate_reg_1[3180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6359]),.i2(intermediate_reg_0[6358]),.o(intermediate_reg_1[3179]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6357]),.i2(intermediate_reg_0[6356]),.o(intermediate_reg_1[3178]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6355]),.i2(intermediate_reg_0[6354]),.o(intermediate_reg_1[3177]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6353]),.i2(intermediate_reg_0[6352]),.o(intermediate_reg_1[3176])); 
xor_module xor_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6351]),.i2(intermediate_reg_0[6350]),.o(intermediate_reg_1[3175])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6349]),.i2(intermediate_reg_0[6348]),.o(intermediate_reg_1[3174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6347]),.i2(intermediate_reg_0[6346]),.o(intermediate_reg_1[3173]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6345]),.i2(intermediate_reg_0[6344]),.o(intermediate_reg_1[3172])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6343]),.i2(intermediate_reg_0[6342]),.o(intermediate_reg_1[3171]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6341]),.i2(intermediate_reg_0[6340]),.o(intermediate_reg_1[3170])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6339]),.i2(intermediate_reg_0[6338]),.o(intermediate_reg_1[3169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6337]),.i2(intermediate_reg_0[6336]),.o(intermediate_reg_1[3168]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6335]),.i2(intermediate_reg_0[6334]),.o(intermediate_reg_1[3167])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6333]),.i2(intermediate_reg_0[6332]),.o(intermediate_reg_1[3166])); 
xor_module xor_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6331]),.i2(intermediate_reg_0[6330]),.o(intermediate_reg_1[3165])); 
mux_module mux_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6329]),.i2(intermediate_reg_0[6328]),.o(intermediate_reg_1[3164]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6327]),.i2(intermediate_reg_0[6326]),.o(intermediate_reg_1[3163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6325]),.i2(intermediate_reg_0[6324]),.o(intermediate_reg_1[3162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6323]),.i2(intermediate_reg_0[6322]),.o(intermediate_reg_1[3161]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6321]),.i2(intermediate_reg_0[6320]),.o(intermediate_reg_1[3160])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6319]),.i2(intermediate_reg_0[6318]),.o(intermediate_reg_1[3159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6317]),.i2(intermediate_reg_0[6316]),.o(intermediate_reg_1[3158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6315]),.i2(intermediate_reg_0[6314]),.o(intermediate_reg_1[3157]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6313]),.i2(intermediate_reg_0[6312]),.o(intermediate_reg_1[3156])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6311]),.i2(intermediate_reg_0[6310]),.o(intermediate_reg_1[3155])); 
mux_module mux_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6309]),.i2(intermediate_reg_0[6308]),.o(intermediate_reg_1[3154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6307]),.i2(intermediate_reg_0[6306]),.o(intermediate_reg_1[3153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6305]),.i2(intermediate_reg_0[6304]),.o(intermediate_reg_1[3152]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6303]),.i2(intermediate_reg_0[6302]),.o(intermediate_reg_1[3151])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6301]),.i2(intermediate_reg_0[6300]),.o(intermediate_reg_1[3150])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6299]),.i2(intermediate_reg_0[6298]),.o(intermediate_reg_1[3149]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6297]),.i2(intermediate_reg_0[6296]),.o(intermediate_reg_1[3148])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6295]),.i2(intermediate_reg_0[6294]),.o(intermediate_reg_1[3147]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6293]),.i2(intermediate_reg_0[6292]),.o(intermediate_reg_1[3146])); 
mux_module mux_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6291]),.i2(intermediate_reg_0[6290]),.o(intermediate_reg_1[3145]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6289]),.i2(intermediate_reg_0[6288]),.o(intermediate_reg_1[3144])); 
xor_module xor_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6287]),.i2(intermediate_reg_0[6286]),.o(intermediate_reg_1[3143])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6285]),.i2(intermediate_reg_0[6284]),.o(intermediate_reg_1[3142]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6283]),.i2(intermediate_reg_0[6282]),.o(intermediate_reg_1[3141]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6281]),.i2(intermediate_reg_0[6280]),.o(intermediate_reg_1[3140])); 
mux_module mux_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6279]),.i2(intermediate_reg_0[6278]),.o(intermediate_reg_1[3139]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6277]),.i2(intermediate_reg_0[6276]),.o(intermediate_reg_1[3138])); 
mux_module mux_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6275]),.i2(intermediate_reg_0[6274]),.o(intermediate_reg_1[3137]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6273]),.i2(intermediate_reg_0[6272]),.o(intermediate_reg_1[3136])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6271]),.i2(intermediate_reg_0[6270]),.o(intermediate_reg_1[3135]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6269]),.i2(intermediate_reg_0[6268]),.o(intermediate_reg_1[3134])); 
xor_module xor_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6267]),.i2(intermediate_reg_0[6266]),.o(intermediate_reg_1[3133])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6265]),.i2(intermediate_reg_0[6264]),.o(intermediate_reg_1[3132]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6263]),.i2(intermediate_reg_0[6262]),.o(intermediate_reg_1[3131])); 
xor_module xor_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6261]),.i2(intermediate_reg_0[6260]),.o(intermediate_reg_1[3130])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6259]),.i2(intermediate_reg_0[6258]),.o(intermediate_reg_1[3129]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6257]),.i2(intermediate_reg_0[6256]),.o(intermediate_reg_1[3128]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6255]),.i2(intermediate_reg_0[6254]),.o(intermediate_reg_1[3127])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6253]),.i2(intermediate_reg_0[6252]),.o(intermediate_reg_1[3126]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6251]),.i2(intermediate_reg_0[6250]),.o(intermediate_reg_1[3125])); 
xor_module xor_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6249]),.i2(intermediate_reg_0[6248]),.o(intermediate_reg_1[3124])); 
mux_module mux_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6247]),.i2(intermediate_reg_0[6246]),.o(intermediate_reg_1[3123]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6245]),.i2(intermediate_reg_0[6244]),.o(intermediate_reg_1[3122])); 
xor_module xor_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6243]),.i2(intermediate_reg_0[6242]),.o(intermediate_reg_1[3121])); 
mux_module mux_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6241]),.i2(intermediate_reg_0[6240]),.o(intermediate_reg_1[3120]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6239]),.i2(intermediate_reg_0[6238]),.o(intermediate_reg_1[3119])); 
xor_module xor_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6237]),.i2(intermediate_reg_0[6236]),.o(intermediate_reg_1[3118])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6235]),.i2(intermediate_reg_0[6234]),.o(intermediate_reg_1[3117])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6233]),.i2(intermediate_reg_0[6232]),.o(intermediate_reg_1[3116]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6231]),.i2(intermediate_reg_0[6230]),.o(intermediate_reg_1[3115])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6229]),.i2(intermediate_reg_0[6228]),.o(intermediate_reg_1[3114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6227]),.i2(intermediate_reg_0[6226]),.o(intermediate_reg_1[3113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6225]),.i2(intermediate_reg_0[6224]),.o(intermediate_reg_1[3112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6223]),.i2(intermediate_reg_0[6222]),.o(intermediate_reg_1[3111]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6221]),.i2(intermediate_reg_0[6220]),.o(intermediate_reg_1[3110]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6219]),.i2(intermediate_reg_0[6218]),.o(intermediate_reg_1[3109])); 
mux_module mux_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6217]),.i2(intermediate_reg_0[6216]),.o(intermediate_reg_1[3108]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6215]),.i2(intermediate_reg_0[6214]),.o(intermediate_reg_1[3107])); 
xor_module xor_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6213]),.i2(intermediate_reg_0[6212]),.o(intermediate_reg_1[3106])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6211]),.i2(intermediate_reg_0[6210]),.o(intermediate_reg_1[3105]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6209]),.i2(intermediate_reg_0[6208]),.o(intermediate_reg_1[3104]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6207]),.i2(intermediate_reg_0[6206]),.o(intermediate_reg_1[3103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6205]),.i2(intermediate_reg_0[6204]),.o(intermediate_reg_1[3102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6203]),.i2(intermediate_reg_0[6202]),.o(intermediate_reg_1[3101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6201]),.i2(intermediate_reg_0[6200]),.o(intermediate_reg_1[3100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6199]),.i2(intermediate_reg_0[6198]),.o(intermediate_reg_1[3099]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6197]),.i2(intermediate_reg_0[6196]),.o(intermediate_reg_1[3098]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6195]),.i2(intermediate_reg_0[6194]),.o(intermediate_reg_1[3097])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6193]),.i2(intermediate_reg_0[6192]),.o(intermediate_reg_1[3096]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6191]),.i2(intermediate_reg_0[6190]),.o(intermediate_reg_1[3095])); 
xor_module xor_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6189]),.i2(intermediate_reg_0[6188]),.o(intermediate_reg_1[3094])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6187]),.i2(intermediate_reg_0[6186]),.o(intermediate_reg_1[3093]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6185]),.i2(intermediate_reg_0[6184]),.o(intermediate_reg_1[3092])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6183]),.i2(intermediate_reg_0[6182]),.o(intermediate_reg_1[3091]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6181]),.i2(intermediate_reg_0[6180]),.o(intermediate_reg_1[3090])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6179]),.i2(intermediate_reg_0[6178]),.o(intermediate_reg_1[3089]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6177]),.i2(intermediate_reg_0[6176]),.o(intermediate_reg_1[3088]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6175]),.i2(intermediate_reg_0[6174]),.o(intermediate_reg_1[3087]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6173]),.i2(intermediate_reg_0[6172]),.o(intermediate_reg_1[3086])); 
xor_module xor_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6171]),.i2(intermediate_reg_0[6170]),.o(intermediate_reg_1[3085])); 
xor_module xor_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6169]),.i2(intermediate_reg_0[6168]),.o(intermediate_reg_1[3084])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6167]),.i2(intermediate_reg_0[6166]),.o(intermediate_reg_1[3083]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6165]),.i2(intermediate_reg_0[6164]),.o(intermediate_reg_1[3082])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6163]),.i2(intermediate_reg_0[6162]),.o(intermediate_reg_1[3081])); 
xor_module xor_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6161]),.i2(intermediate_reg_0[6160]),.o(intermediate_reg_1[3080])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6159]),.i2(intermediate_reg_0[6158]),.o(intermediate_reg_1[3079]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6157]),.i2(intermediate_reg_0[6156]),.o(intermediate_reg_1[3078])); 
mux_module mux_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6155]),.i2(intermediate_reg_0[6154]),.o(intermediate_reg_1[3077]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6153]),.i2(intermediate_reg_0[6152]),.o(intermediate_reg_1[3076]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6151]),.i2(intermediate_reg_0[6150]),.o(intermediate_reg_1[3075]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6149]),.i2(intermediate_reg_0[6148]),.o(intermediate_reg_1[3074])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6147]),.i2(intermediate_reg_0[6146]),.o(intermediate_reg_1[3073])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6145]),.i2(intermediate_reg_0[6144]),.o(intermediate_reg_1[3072])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6143]),.i2(intermediate_reg_0[6142]),.o(intermediate_reg_1[3071])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6141]),.i2(intermediate_reg_0[6140]),.o(intermediate_reg_1[3070])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6139]),.i2(intermediate_reg_0[6138]),.o(intermediate_reg_1[3069])); 
xor_module xor_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6137]),.i2(intermediate_reg_0[6136]),.o(intermediate_reg_1[3068])); 
xor_module xor_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6135]),.i2(intermediate_reg_0[6134]),.o(intermediate_reg_1[3067])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6133]),.i2(intermediate_reg_0[6132]),.o(intermediate_reg_1[3066]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6131]),.i2(intermediate_reg_0[6130]),.o(intermediate_reg_1[3065]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6129]),.i2(intermediate_reg_0[6128]),.o(intermediate_reg_1[3064])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6127]),.i2(intermediate_reg_0[6126]),.o(intermediate_reg_1[3063]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6125]),.i2(intermediate_reg_0[6124]),.o(intermediate_reg_1[3062]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6123]),.i2(intermediate_reg_0[6122]),.o(intermediate_reg_1[3061])); 
mux_module mux_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6121]),.i2(intermediate_reg_0[6120]),.o(intermediate_reg_1[3060]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6119]),.i2(intermediate_reg_0[6118]),.o(intermediate_reg_1[3059])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6117]),.i2(intermediate_reg_0[6116]),.o(intermediate_reg_1[3058]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6115]),.i2(intermediate_reg_0[6114]),.o(intermediate_reg_1[3057]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6113]),.i2(intermediate_reg_0[6112]),.o(intermediate_reg_1[3056]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6111]),.i2(intermediate_reg_0[6110]),.o(intermediate_reg_1[3055])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6109]),.i2(intermediate_reg_0[6108]),.o(intermediate_reg_1[3054])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6107]),.i2(intermediate_reg_0[6106]),.o(intermediate_reg_1[3053]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6105]),.i2(intermediate_reg_0[6104]),.o(intermediate_reg_1[3052])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6103]),.i2(intermediate_reg_0[6102]),.o(intermediate_reg_1[3051]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6101]),.i2(intermediate_reg_0[6100]),.o(intermediate_reg_1[3050])); 
xor_module xor_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6099]),.i2(intermediate_reg_0[6098]),.o(intermediate_reg_1[3049])); 
xor_module xor_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6097]),.i2(intermediate_reg_0[6096]),.o(intermediate_reg_1[3048])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6095]),.i2(intermediate_reg_0[6094]),.o(intermediate_reg_1[3047])); 
mux_module mux_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6093]),.i2(intermediate_reg_0[6092]),.o(intermediate_reg_1[3046]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6091]),.i2(intermediate_reg_0[6090]),.o(intermediate_reg_1[3045]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6089]),.i2(intermediate_reg_0[6088]),.o(intermediate_reg_1[3044])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6087]),.i2(intermediate_reg_0[6086]),.o(intermediate_reg_1[3043]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6085]),.i2(intermediate_reg_0[6084]),.o(intermediate_reg_1[3042])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6083]),.i2(intermediate_reg_0[6082]),.o(intermediate_reg_1[3041]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6081]),.i2(intermediate_reg_0[6080]),.o(intermediate_reg_1[3040])); 
mux_module mux_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6079]),.i2(intermediate_reg_0[6078]),.o(intermediate_reg_1[3039]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6077]),.i2(intermediate_reg_0[6076]),.o(intermediate_reg_1[3038])); 
xor_module xor_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6075]),.i2(intermediate_reg_0[6074]),.o(intermediate_reg_1[3037])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6073]),.i2(intermediate_reg_0[6072]),.o(intermediate_reg_1[3036]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6071]),.i2(intermediate_reg_0[6070]),.o(intermediate_reg_1[3035]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6069]),.i2(intermediate_reg_0[6068]),.o(intermediate_reg_1[3034]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6067]),.i2(intermediate_reg_0[6066]),.o(intermediate_reg_1[3033]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6065]),.i2(intermediate_reg_0[6064]),.o(intermediate_reg_1[3032]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6063]),.i2(intermediate_reg_0[6062]),.o(intermediate_reg_1[3031])); 
xor_module xor_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6061]),.i2(intermediate_reg_0[6060]),.o(intermediate_reg_1[3030])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6059]),.i2(intermediate_reg_0[6058]),.o(intermediate_reg_1[3029])); 
xor_module xor_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6057]),.i2(intermediate_reg_0[6056]),.o(intermediate_reg_1[3028])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6055]),.i2(intermediate_reg_0[6054]),.o(intermediate_reg_1[3027]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6053]),.i2(intermediate_reg_0[6052]),.o(intermediate_reg_1[3026])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6051]),.i2(intermediate_reg_0[6050]),.o(intermediate_reg_1[3025]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6049]),.i2(intermediate_reg_0[6048]),.o(intermediate_reg_1[3024])); 
xor_module xor_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6047]),.i2(intermediate_reg_0[6046]),.o(intermediate_reg_1[3023])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6045]),.i2(intermediate_reg_0[6044]),.o(intermediate_reg_1[3022]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6043]),.i2(intermediate_reg_0[6042]),.o(intermediate_reg_1[3021]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6041]),.i2(intermediate_reg_0[6040]),.o(intermediate_reg_1[3020])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6039]),.i2(intermediate_reg_0[6038]),.o(intermediate_reg_1[3019]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6037]),.i2(intermediate_reg_0[6036]),.o(intermediate_reg_1[3018]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6035]),.i2(intermediate_reg_0[6034]),.o(intermediate_reg_1[3017])); 
xor_module xor_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6033]),.i2(intermediate_reg_0[6032]),.o(intermediate_reg_1[3016])); 
xor_module xor_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6031]),.i2(intermediate_reg_0[6030]),.o(intermediate_reg_1[3015])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6029]),.i2(intermediate_reg_0[6028]),.o(intermediate_reg_1[3014])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6027]),.i2(intermediate_reg_0[6026]),.o(intermediate_reg_1[3013]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6025]),.i2(intermediate_reg_0[6024]),.o(intermediate_reg_1[3012])); 
xor_module xor_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6023]),.i2(intermediate_reg_0[6022]),.o(intermediate_reg_1[3011])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6021]),.i2(intermediate_reg_0[6020]),.o(intermediate_reg_1[3010])); 
xor_module xor_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6019]),.i2(intermediate_reg_0[6018]),.o(intermediate_reg_1[3009])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6017]),.i2(intermediate_reg_0[6016]),.o(intermediate_reg_1[3008]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6015]),.i2(intermediate_reg_0[6014]),.o(intermediate_reg_1[3007])); 
mux_module mux_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6013]),.i2(intermediate_reg_0[6012]),.o(intermediate_reg_1[3006]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6011]),.i2(intermediate_reg_0[6010]),.o(intermediate_reg_1[3005])); 
mux_module mux_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6009]),.i2(intermediate_reg_0[6008]),.o(intermediate_reg_1[3004]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6007]),.i2(intermediate_reg_0[6006]),.o(intermediate_reg_1[3003]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6005]),.i2(intermediate_reg_0[6004]),.o(intermediate_reg_1[3002])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6003]),.i2(intermediate_reg_0[6002]),.o(intermediate_reg_1[3001]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6001]),.i2(intermediate_reg_0[6000]),.o(intermediate_reg_1[3000]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5999]),.i2(intermediate_reg_0[5998]),.o(intermediate_reg_1[2999]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5997]),.i2(intermediate_reg_0[5996]),.o(intermediate_reg_1[2998]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5995]),.i2(intermediate_reg_0[5994]),.o(intermediate_reg_1[2997]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5993]),.i2(intermediate_reg_0[5992]),.o(intermediate_reg_1[2996]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5991]),.i2(intermediate_reg_0[5990]),.o(intermediate_reg_1[2995]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5989]),.i2(intermediate_reg_0[5988]),.o(intermediate_reg_1[2994])); 
mux_module mux_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5987]),.i2(intermediate_reg_0[5986]),.o(intermediate_reg_1[2993]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5985]),.i2(intermediate_reg_0[5984]),.o(intermediate_reg_1[2992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5983]),.i2(intermediate_reg_0[5982]),.o(intermediate_reg_1[2991]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5981]),.i2(intermediate_reg_0[5980]),.o(intermediate_reg_1[2990])); 
mux_module mux_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5979]),.i2(intermediate_reg_0[5978]),.o(intermediate_reg_1[2989]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5977]),.i2(intermediate_reg_0[5976]),.o(intermediate_reg_1[2988])); 
xor_module xor_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5975]),.i2(intermediate_reg_0[5974]),.o(intermediate_reg_1[2987])); 
xor_module xor_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5973]),.i2(intermediate_reg_0[5972]),.o(intermediate_reg_1[2986])); 
mux_module mux_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5971]),.i2(intermediate_reg_0[5970]),.o(intermediate_reg_1[2985]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5969]),.i2(intermediate_reg_0[5968]),.o(intermediate_reg_1[2984])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5967]),.i2(intermediate_reg_0[5966]),.o(intermediate_reg_1[2983]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5965]),.i2(intermediate_reg_0[5964]),.o(intermediate_reg_1[2982])); 
mux_module mux_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5963]),.i2(intermediate_reg_0[5962]),.o(intermediate_reg_1[2981]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5961]),.i2(intermediate_reg_0[5960]),.o(intermediate_reg_1[2980]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5959]),.i2(intermediate_reg_0[5958]),.o(intermediate_reg_1[2979])); 
mux_module mux_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5957]),.i2(intermediate_reg_0[5956]),.o(intermediate_reg_1[2978]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5955]),.i2(intermediate_reg_0[5954]),.o(intermediate_reg_1[2977])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5953]),.i2(intermediate_reg_0[5952]),.o(intermediate_reg_1[2976]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5951]),.i2(intermediate_reg_0[5950]),.o(intermediate_reg_1[2975])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5949]),.i2(intermediate_reg_0[5948]),.o(intermediate_reg_1[2974]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5947]),.i2(intermediate_reg_0[5946]),.o(intermediate_reg_1[2973])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5945]),.i2(intermediate_reg_0[5944]),.o(intermediate_reg_1[2972]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5943]),.i2(intermediate_reg_0[5942]),.o(intermediate_reg_1[2971])); 
xor_module xor_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5941]),.i2(intermediate_reg_0[5940]),.o(intermediate_reg_1[2970])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5939]),.i2(intermediate_reg_0[5938]),.o(intermediate_reg_1[2969])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5937]),.i2(intermediate_reg_0[5936]),.o(intermediate_reg_1[2968])); 
xor_module xor_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5935]),.i2(intermediate_reg_0[5934]),.o(intermediate_reg_1[2967])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5933]),.i2(intermediate_reg_0[5932]),.o(intermediate_reg_1[2966]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5931]),.i2(intermediate_reg_0[5930]),.o(intermediate_reg_1[2965])); 
mux_module mux_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5929]),.i2(intermediate_reg_0[5928]),.o(intermediate_reg_1[2964]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5927]),.i2(intermediate_reg_0[5926]),.o(intermediate_reg_1[2963])); 
xor_module xor_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5925]),.i2(intermediate_reg_0[5924]),.o(intermediate_reg_1[2962])); 
mux_module mux_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5923]),.i2(intermediate_reg_0[5922]),.o(intermediate_reg_1[2961]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5921]),.i2(intermediate_reg_0[5920]),.o(intermediate_reg_1[2960])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5919]),.i2(intermediate_reg_0[5918]),.o(intermediate_reg_1[2959]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5917]),.i2(intermediate_reg_0[5916]),.o(intermediate_reg_1[2958])); 
xor_module xor_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5915]),.i2(intermediate_reg_0[5914]),.o(intermediate_reg_1[2957])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5913]),.i2(intermediate_reg_0[5912]),.o(intermediate_reg_1[2956])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5911]),.i2(intermediate_reg_0[5910]),.o(intermediate_reg_1[2955]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5909]),.i2(intermediate_reg_0[5908]),.o(intermediate_reg_1[2954]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5907]),.i2(intermediate_reg_0[5906]),.o(intermediate_reg_1[2953])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5905]),.i2(intermediate_reg_0[5904]),.o(intermediate_reg_1[2952])); 
mux_module mux_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5903]),.i2(intermediate_reg_0[5902]),.o(intermediate_reg_1[2951]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5901]),.i2(intermediate_reg_0[5900]),.o(intermediate_reg_1[2950])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5899]),.i2(intermediate_reg_0[5898]),.o(intermediate_reg_1[2949]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5897]),.i2(intermediate_reg_0[5896]),.o(intermediate_reg_1[2948]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5895]),.i2(intermediate_reg_0[5894]),.o(intermediate_reg_1[2947])); 
xor_module xor_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5893]),.i2(intermediate_reg_0[5892]),.o(intermediate_reg_1[2946])); 
xor_module xor_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5891]),.i2(intermediate_reg_0[5890]),.o(intermediate_reg_1[2945])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5889]),.i2(intermediate_reg_0[5888]),.o(intermediate_reg_1[2944])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5887]),.i2(intermediate_reg_0[5886]),.o(intermediate_reg_1[2943])); 
xor_module xor_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5885]),.i2(intermediate_reg_0[5884]),.o(intermediate_reg_1[2942])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5883]),.i2(intermediate_reg_0[5882]),.o(intermediate_reg_1[2941])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5881]),.i2(intermediate_reg_0[5880]),.o(intermediate_reg_1[2940]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5879]),.i2(intermediate_reg_0[5878]),.o(intermediate_reg_1[2939]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5877]),.i2(intermediate_reg_0[5876]),.o(intermediate_reg_1[2938])); 
mux_module mux_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5875]),.i2(intermediate_reg_0[5874]),.o(intermediate_reg_1[2937]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5873]),.i2(intermediate_reg_0[5872]),.o(intermediate_reg_1[2936]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5871]),.i2(intermediate_reg_0[5870]),.o(intermediate_reg_1[2935])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5869]),.i2(intermediate_reg_0[5868]),.o(intermediate_reg_1[2934])); 
mux_module mux_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5867]),.i2(intermediate_reg_0[5866]),.o(intermediate_reg_1[2933]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5865]),.i2(intermediate_reg_0[5864]),.o(intermediate_reg_1[2932]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5863]),.i2(intermediate_reg_0[5862]),.o(intermediate_reg_1[2931])); 
xor_module xor_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5861]),.i2(intermediate_reg_0[5860]),.o(intermediate_reg_1[2930])); 
xor_module xor_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5859]),.i2(intermediate_reg_0[5858]),.o(intermediate_reg_1[2929])); 
xor_module xor_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5857]),.i2(intermediate_reg_0[5856]),.o(intermediate_reg_1[2928])); 
xor_module xor_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5855]),.i2(intermediate_reg_0[5854]),.o(intermediate_reg_1[2927])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5853]),.i2(intermediate_reg_0[5852]),.o(intermediate_reg_1[2926]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5851]),.i2(intermediate_reg_0[5850]),.o(intermediate_reg_1[2925])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5849]),.i2(intermediate_reg_0[5848]),.o(intermediate_reg_1[2924]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5847]),.i2(intermediate_reg_0[5846]),.o(intermediate_reg_1[2923])); 
xor_module xor_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5845]),.i2(intermediate_reg_0[5844]),.o(intermediate_reg_1[2922])); 
mux_module mux_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5843]),.i2(intermediate_reg_0[5842]),.o(intermediate_reg_1[2921]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5841]),.i2(intermediate_reg_0[5840]),.o(intermediate_reg_1[2920])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5839]),.i2(intermediate_reg_0[5838]),.o(intermediate_reg_1[2919])); 
xor_module xor_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5837]),.i2(intermediate_reg_0[5836]),.o(intermediate_reg_1[2918])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5835]),.i2(intermediate_reg_0[5834]),.o(intermediate_reg_1[2917]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5833]),.i2(intermediate_reg_0[5832]),.o(intermediate_reg_1[2916]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5831]),.i2(intermediate_reg_0[5830]),.o(intermediate_reg_1[2915])); 
mux_module mux_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5829]),.i2(intermediate_reg_0[5828]),.o(intermediate_reg_1[2914]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5827]),.i2(intermediate_reg_0[5826]),.o(intermediate_reg_1[2913])); 
xor_module xor_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5825]),.i2(intermediate_reg_0[5824]),.o(intermediate_reg_1[2912])); 
mux_module mux_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5823]),.i2(intermediate_reg_0[5822]),.o(intermediate_reg_1[2911]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5821]),.i2(intermediate_reg_0[5820]),.o(intermediate_reg_1[2910]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5819]),.i2(intermediate_reg_0[5818]),.o(intermediate_reg_1[2909])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5817]),.i2(intermediate_reg_0[5816]),.o(intermediate_reg_1[2908]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5815]),.i2(intermediate_reg_0[5814]),.o(intermediate_reg_1[2907])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5813]),.i2(intermediate_reg_0[5812]),.o(intermediate_reg_1[2906])); 
mux_module mux_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5811]),.i2(intermediate_reg_0[5810]),.o(intermediate_reg_1[2905]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5809]),.i2(intermediate_reg_0[5808]),.o(intermediate_reg_1[2904])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5807]),.i2(intermediate_reg_0[5806]),.o(intermediate_reg_1[2903]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5805]),.i2(intermediate_reg_0[5804]),.o(intermediate_reg_1[2902])); 
xor_module xor_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5803]),.i2(intermediate_reg_0[5802]),.o(intermediate_reg_1[2901])); 
xor_module xor_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5801]),.i2(intermediate_reg_0[5800]),.o(intermediate_reg_1[2900])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5799]),.i2(intermediate_reg_0[5798]),.o(intermediate_reg_1[2899])); 
xor_module xor_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5797]),.i2(intermediate_reg_0[5796]),.o(intermediate_reg_1[2898])); 
xor_module xor_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5795]),.i2(intermediate_reg_0[5794]),.o(intermediate_reg_1[2897])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5793]),.i2(intermediate_reg_0[5792]),.o(intermediate_reg_1[2896]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5791]),.i2(intermediate_reg_0[5790]),.o(intermediate_reg_1[2895])); 
mux_module mux_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5789]),.i2(intermediate_reg_0[5788]),.o(intermediate_reg_1[2894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5787]),.i2(intermediate_reg_0[5786]),.o(intermediate_reg_1[2893]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5785]),.i2(intermediate_reg_0[5784]),.o(intermediate_reg_1[2892]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5783]),.i2(intermediate_reg_0[5782]),.o(intermediate_reg_1[2891]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5781]),.i2(intermediate_reg_0[5780]),.o(intermediate_reg_1[2890]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5779]),.i2(intermediate_reg_0[5778]),.o(intermediate_reg_1[2889])); 
xor_module xor_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5777]),.i2(intermediate_reg_0[5776]),.o(intermediate_reg_1[2888])); 
mux_module mux_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5775]),.i2(intermediate_reg_0[5774]),.o(intermediate_reg_1[2887]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5773]),.i2(intermediate_reg_0[5772]),.o(intermediate_reg_1[2886])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5771]),.i2(intermediate_reg_0[5770]),.o(intermediate_reg_1[2885])); 
xor_module xor_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5769]),.i2(intermediate_reg_0[5768]),.o(intermediate_reg_1[2884])); 
xor_module xor_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5767]),.i2(intermediate_reg_0[5766]),.o(intermediate_reg_1[2883])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5765]),.i2(intermediate_reg_0[5764]),.o(intermediate_reg_1[2882])); 
mux_module mux_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5763]),.i2(intermediate_reg_0[5762]),.o(intermediate_reg_1[2881]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5761]),.i2(intermediate_reg_0[5760]),.o(intermediate_reg_1[2880]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5759]),.i2(intermediate_reg_0[5758]),.o(intermediate_reg_1[2879]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5757]),.i2(intermediate_reg_0[5756]),.o(intermediate_reg_1[2878]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5755]),.i2(intermediate_reg_0[5754]),.o(intermediate_reg_1[2877])); 
mux_module mux_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5753]),.i2(intermediate_reg_0[5752]),.o(intermediate_reg_1[2876]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5751]),.i2(intermediate_reg_0[5750]),.o(intermediate_reg_1[2875])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5749]),.i2(intermediate_reg_0[5748]),.o(intermediate_reg_1[2874]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5747]),.i2(intermediate_reg_0[5746]),.o(intermediate_reg_1[2873]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5745]),.i2(intermediate_reg_0[5744]),.o(intermediate_reg_1[2872]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5743]),.i2(intermediate_reg_0[5742]),.o(intermediate_reg_1[2871])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5741]),.i2(intermediate_reg_0[5740]),.o(intermediate_reg_1[2870]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5739]),.i2(intermediate_reg_0[5738]),.o(intermediate_reg_1[2869])); 
xor_module xor_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5737]),.i2(intermediate_reg_0[5736]),.o(intermediate_reg_1[2868])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5735]),.i2(intermediate_reg_0[5734]),.o(intermediate_reg_1[2867])); 
xor_module xor_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5733]),.i2(intermediate_reg_0[5732]),.o(intermediate_reg_1[2866])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5731]),.i2(intermediate_reg_0[5730]),.o(intermediate_reg_1[2865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5729]),.i2(intermediate_reg_0[5728]),.o(intermediate_reg_1[2864]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5727]),.i2(intermediate_reg_0[5726]),.o(intermediate_reg_1[2863])); 
mux_module mux_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5725]),.i2(intermediate_reg_0[5724]),.o(intermediate_reg_1[2862]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5723]),.i2(intermediate_reg_0[5722]),.o(intermediate_reg_1[2861]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5721]),.i2(intermediate_reg_0[5720]),.o(intermediate_reg_1[2860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5719]),.i2(intermediate_reg_0[5718]),.o(intermediate_reg_1[2859]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5717]),.i2(intermediate_reg_0[5716]),.o(intermediate_reg_1[2858])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5715]),.i2(intermediate_reg_0[5714]),.o(intermediate_reg_1[2857]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5713]),.i2(intermediate_reg_0[5712]),.o(intermediate_reg_1[2856])); 
xor_module xor_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5711]),.i2(intermediate_reg_0[5710]),.o(intermediate_reg_1[2855])); 
xor_module xor_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5709]),.i2(intermediate_reg_0[5708]),.o(intermediate_reg_1[2854])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5707]),.i2(intermediate_reg_0[5706]),.o(intermediate_reg_1[2853])); 
mux_module mux_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5705]),.i2(intermediate_reg_0[5704]),.o(intermediate_reg_1[2852]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5703]),.i2(intermediate_reg_0[5702]),.o(intermediate_reg_1[2851])); 
mux_module mux_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5701]),.i2(intermediate_reg_0[5700]),.o(intermediate_reg_1[2850]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5699]),.i2(intermediate_reg_0[5698]),.o(intermediate_reg_1[2849])); 
xor_module xor_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5697]),.i2(intermediate_reg_0[5696]),.o(intermediate_reg_1[2848])); 
xor_module xor_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5695]),.i2(intermediate_reg_0[5694]),.o(intermediate_reg_1[2847])); 
mux_module mux_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5693]),.i2(intermediate_reg_0[5692]),.o(intermediate_reg_1[2846]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5691]),.i2(intermediate_reg_0[5690]),.o(intermediate_reg_1[2845]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5689]),.i2(intermediate_reg_0[5688]),.o(intermediate_reg_1[2844]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5687]),.i2(intermediate_reg_0[5686]),.o(intermediate_reg_1[2843]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5685]),.i2(intermediate_reg_0[5684]),.o(intermediate_reg_1[2842]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5683]),.i2(intermediate_reg_0[5682]),.o(intermediate_reg_1[2841])); 
xor_module xor_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5681]),.i2(intermediate_reg_0[5680]),.o(intermediate_reg_1[2840])); 
mux_module mux_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5679]),.i2(intermediate_reg_0[5678]),.o(intermediate_reg_1[2839]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5677]),.i2(intermediate_reg_0[5676]),.o(intermediate_reg_1[2838])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5675]),.i2(intermediate_reg_0[5674]),.o(intermediate_reg_1[2837]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5673]),.i2(intermediate_reg_0[5672]),.o(intermediate_reg_1[2836])); 
mux_module mux_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5671]),.i2(intermediate_reg_0[5670]),.o(intermediate_reg_1[2835]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5669]),.i2(intermediate_reg_0[5668]),.o(intermediate_reg_1[2834]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5667]),.i2(intermediate_reg_0[5666]),.o(intermediate_reg_1[2833])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5665]),.i2(intermediate_reg_0[5664]),.o(intermediate_reg_1[2832])); 
xor_module xor_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5663]),.i2(intermediate_reg_0[5662]),.o(intermediate_reg_1[2831])); 
mux_module mux_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5661]),.i2(intermediate_reg_0[5660]),.o(intermediate_reg_1[2830]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5659]),.i2(intermediate_reg_0[5658]),.o(intermediate_reg_1[2829])); 
xor_module xor_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5657]),.i2(intermediate_reg_0[5656]),.o(intermediate_reg_1[2828])); 
xor_module xor_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5655]),.i2(intermediate_reg_0[5654]),.o(intermediate_reg_1[2827])); 
xor_module xor_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5653]),.i2(intermediate_reg_0[5652]),.o(intermediate_reg_1[2826])); 
mux_module mux_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5651]),.i2(intermediate_reg_0[5650]),.o(intermediate_reg_1[2825]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5649]),.i2(intermediate_reg_0[5648]),.o(intermediate_reg_1[2824]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5647]),.i2(intermediate_reg_0[5646]),.o(intermediate_reg_1[2823])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5645]),.i2(intermediate_reg_0[5644]),.o(intermediate_reg_1[2822]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5643]),.i2(intermediate_reg_0[5642]),.o(intermediate_reg_1[2821])); 
mux_module mux_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5641]),.i2(intermediate_reg_0[5640]),.o(intermediate_reg_1[2820]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5639]),.i2(intermediate_reg_0[5638]),.o(intermediate_reg_1[2819])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5637]),.i2(intermediate_reg_0[5636]),.o(intermediate_reg_1[2818]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5635]),.i2(intermediate_reg_0[5634]),.o(intermediate_reg_1[2817])); 
xor_module xor_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5633]),.i2(intermediate_reg_0[5632]),.o(intermediate_reg_1[2816])); 
mux_module mux_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5631]),.i2(intermediate_reg_0[5630]),.o(intermediate_reg_1[2815]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5629]),.i2(intermediate_reg_0[5628]),.o(intermediate_reg_1[2814]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5627]),.i2(intermediate_reg_0[5626]),.o(intermediate_reg_1[2813]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5625]),.i2(intermediate_reg_0[5624]),.o(intermediate_reg_1[2812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5623]),.i2(intermediate_reg_0[5622]),.o(intermediate_reg_1[2811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5621]),.i2(intermediate_reg_0[5620]),.o(intermediate_reg_1[2810]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5619]),.i2(intermediate_reg_0[5618]),.o(intermediate_reg_1[2809])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5617]),.i2(intermediate_reg_0[5616]),.o(intermediate_reg_1[2808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5615]),.i2(intermediate_reg_0[5614]),.o(intermediate_reg_1[2807]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5613]),.i2(intermediate_reg_0[5612]),.o(intermediate_reg_1[2806])); 
mux_module mux_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5611]),.i2(intermediate_reg_0[5610]),.o(intermediate_reg_1[2805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5609]),.i2(intermediate_reg_0[5608]),.o(intermediate_reg_1[2804]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5607]),.i2(intermediate_reg_0[5606]),.o(intermediate_reg_1[2803]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5605]),.i2(intermediate_reg_0[5604]),.o(intermediate_reg_1[2802]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5603]),.i2(intermediate_reg_0[5602]),.o(intermediate_reg_1[2801]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5601]),.i2(intermediate_reg_0[5600]),.o(intermediate_reg_1[2800])); 
xor_module xor_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5599]),.i2(intermediate_reg_0[5598]),.o(intermediate_reg_1[2799])); 
mux_module mux_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5597]),.i2(intermediate_reg_0[5596]),.o(intermediate_reg_1[2798]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5595]),.i2(intermediate_reg_0[5594]),.o(intermediate_reg_1[2797]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5593]),.i2(intermediate_reg_0[5592]),.o(intermediate_reg_1[2796])); 
xor_module xor_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5591]),.i2(intermediate_reg_0[5590]),.o(intermediate_reg_1[2795])); 
mux_module mux_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5589]),.i2(intermediate_reg_0[5588]),.o(intermediate_reg_1[2794]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5587]),.i2(intermediate_reg_0[5586]),.o(intermediate_reg_1[2793])); 
mux_module mux_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5585]),.i2(intermediate_reg_0[5584]),.o(intermediate_reg_1[2792]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5583]),.i2(intermediate_reg_0[5582]),.o(intermediate_reg_1[2791]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5581]),.i2(intermediate_reg_0[5580]),.o(intermediate_reg_1[2790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5579]),.i2(intermediate_reg_0[5578]),.o(intermediate_reg_1[2789]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5577]),.i2(intermediate_reg_0[5576]),.o(intermediate_reg_1[2788])); 
mux_module mux_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5575]),.i2(intermediate_reg_0[5574]),.o(intermediate_reg_1[2787]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5573]),.i2(intermediate_reg_0[5572]),.o(intermediate_reg_1[2786]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5571]),.i2(intermediate_reg_0[5570]),.o(intermediate_reg_1[2785])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5569]),.i2(intermediate_reg_0[5568]),.o(intermediate_reg_1[2784])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5567]),.i2(intermediate_reg_0[5566]),.o(intermediate_reg_1[2783]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5565]),.i2(intermediate_reg_0[5564]),.o(intermediate_reg_1[2782]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5563]),.i2(intermediate_reg_0[5562]),.o(intermediate_reg_1[2781])); 
mux_module mux_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5561]),.i2(intermediate_reg_0[5560]),.o(intermediate_reg_1[2780]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5559]),.i2(intermediate_reg_0[5558]),.o(intermediate_reg_1[2779])); 
xor_module xor_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5557]),.i2(intermediate_reg_0[5556]),.o(intermediate_reg_1[2778])); 
xor_module xor_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5555]),.i2(intermediate_reg_0[5554]),.o(intermediate_reg_1[2777])); 
xor_module xor_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5553]),.i2(intermediate_reg_0[5552]),.o(intermediate_reg_1[2776])); 
xor_module xor_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5551]),.i2(intermediate_reg_0[5550]),.o(intermediate_reg_1[2775])); 
xor_module xor_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5549]),.i2(intermediate_reg_0[5548]),.o(intermediate_reg_1[2774])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5547]),.i2(intermediate_reg_0[5546]),.o(intermediate_reg_1[2773]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5545]),.i2(intermediate_reg_0[5544]),.o(intermediate_reg_1[2772])); 
mux_module mux_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5543]),.i2(intermediate_reg_0[5542]),.o(intermediate_reg_1[2771]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5541]),.i2(intermediate_reg_0[5540]),.o(intermediate_reg_1[2770])); 
mux_module mux_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5539]),.i2(intermediate_reg_0[5538]),.o(intermediate_reg_1[2769]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5537]),.i2(intermediate_reg_0[5536]),.o(intermediate_reg_1[2768])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5535]),.i2(intermediate_reg_0[5534]),.o(intermediate_reg_1[2767]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5533]),.i2(intermediate_reg_0[5532]),.o(intermediate_reg_1[2766]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5531]),.i2(intermediate_reg_0[5530]),.o(intermediate_reg_1[2765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5529]),.i2(intermediate_reg_0[5528]),.o(intermediate_reg_1[2764]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5527]),.i2(intermediate_reg_0[5526]),.o(intermediate_reg_1[2763]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5525]),.i2(intermediate_reg_0[5524]),.o(intermediate_reg_1[2762])); 
xor_module xor_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5523]),.i2(intermediate_reg_0[5522]),.o(intermediate_reg_1[2761])); 
xor_module xor_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5521]),.i2(intermediate_reg_0[5520]),.o(intermediate_reg_1[2760])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5519]),.i2(intermediate_reg_0[5518]),.o(intermediate_reg_1[2759]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5517]),.i2(intermediate_reg_0[5516]),.o(intermediate_reg_1[2758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5515]),.i2(intermediate_reg_0[5514]),.o(intermediate_reg_1[2757]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5513]),.i2(intermediate_reg_0[5512]),.o(intermediate_reg_1[2756])); 
mux_module mux_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5511]),.i2(intermediate_reg_0[5510]),.o(intermediate_reg_1[2755]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5509]),.i2(intermediate_reg_0[5508]),.o(intermediate_reg_1[2754])); 
xor_module xor_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5507]),.i2(intermediate_reg_0[5506]),.o(intermediate_reg_1[2753])); 
mux_module mux_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5505]),.i2(intermediate_reg_0[5504]),.o(intermediate_reg_1[2752]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5503]),.i2(intermediate_reg_0[5502]),.o(intermediate_reg_1[2751])); 
xor_module xor_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5501]),.i2(intermediate_reg_0[5500]),.o(intermediate_reg_1[2750])); 
xor_module xor_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5499]),.i2(intermediate_reg_0[5498]),.o(intermediate_reg_1[2749])); 
xor_module xor_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5497]),.i2(intermediate_reg_0[5496]),.o(intermediate_reg_1[2748])); 
xor_module xor_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5495]),.i2(intermediate_reg_0[5494]),.o(intermediate_reg_1[2747])); 
xor_module xor_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5493]),.i2(intermediate_reg_0[5492]),.o(intermediate_reg_1[2746])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5491]),.i2(intermediate_reg_0[5490]),.o(intermediate_reg_1[2745])); 
mux_module mux_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5489]),.i2(intermediate_reg_0[5488]),.o(intermediate_reg_1[2744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5487]),.i2(intermediate_reg_0[5486]),.o(intermediate_reg_1[2743]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5485]),.i2(intermediate_reg_0[5484]),.o(intermediate_reg_1[2742])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5483]),.i2(intermediate_reg_0[5482]),.o(intermediate_reg_1[2741]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5481]),.i2(intermediate_reg_0[5480]),.o(intermediate_reg_1[2740]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5479]),.i2(intermediate_reg_0[5478]),.o(intermediate_reg_1[2739])); 
xor_module xor_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5477]),.i2(intermediate_reg_0[5476]),.o(intermediate_reg_1[2738])); 
xor_module xor_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5475]),.i2(intermediate_reg_0[5474]),.o(intermediate_reg_1[2737])); 
xor_module xor_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5473]),.i2(intermediate_reg_0[5472]),.o(intermediate_reg_1[2736])); 
mux_module mux_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5471]),.i2(intermediate_reg_0[5470]),.o(intermediate_reg_1[2735]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5469]),.i2(intermediate_reg_0[5468]),.o(intermediate_reg_1[2734])); 
xor_module xor_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5467]),.i2(intermediate_reg_0[5466]),.o(intermediate_reg_1[2733])); 
mux_module mux_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5465]),.i2(intermediate_reg_0[5464]),.o(intermediate_reg_1[2732]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5463]),.i2(intermediate_reg_0[5462]),.o(intermediate_reg_1[2731]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5461]),.i2(intermediate_reg_0[5460]),.o(intermediate_reg_1[2730]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5459]),.i2(intermediate_reg_0[5458]),.o(intermediate_reg_1[2729]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5457]),.i2(intermediate_reg_0[5456]),.o(intermediate_reg_1[2728])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5455]),.i2(intermediate_reg_0[5454]),.o(intermediate_reg_1[2727]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5453]),.i2(intermediate_reg_0[5452]),.o(intermediate_reg_1[2726])); 
xor_module xor_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5451]),.i2(intermediate_reg_0[5450]),.o(intermediate_reg_1[2725])); 
mux_module mux_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5449]),.i2(intermediate_reg_0[5448]),.o(intermediate_reg_1[2724]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5447]),.i2(intermediate_reg_0[5446]),.o(intermediate_reg_1[2723])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5445]),.i2(intermediate_reg_0[5444]),.o(intermediate_reg_1[2722]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5443]),.i2(intermediate_reg_0[5442]),.o(intermediate_reg_1[2721])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5441]),.i2(intermediate_reg_0[5440]),.o(intermediate_reg_1[2720]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5439]),.i2(intermediate_reg_0[5438]),.o(intermediate_reg_1[2719]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5437]),.i2(intermediate_reg_0[5436]),.o(intermediate_reg_1[2718])); 
mux_module mux_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5435]),.i2(intermediate_reg_0[5434]),.o(intermediate_reg_1[2717]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5433]),.i2(intermediate_reg_0[5432]),.o(intermediate_reg_1[2716]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5431]),.i2(intermediate_reg_0[5430]),.o(intermediate_reg_1[2715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5429]),.i2(intermediate_reg_0[5428]),.o(intermediate_reg_1[2714]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5427]),.i2(intermediate_reg_0[5426]),.o(intermediate_reg_1[2713]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5425]),.i2(intermediate_reg_0[5424]),.o(intermediate_reg_1[2712])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5423]),.i2(intermediate_reg_0[5422]),.o(intermediate_reg_1[2711]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5421]),.i2(intermediate_reg_0[5420]),.o(intermediate_reg_1[2710])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5419]),.i2(intermediate_reg_0[5418]),.o(intermediate_reg_1[2709]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5417]),.i2(intermediate_reg_0[5416]),.o(intermediate_reg_1[2708])); 
xor_module xor_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5415]),.i2(intermediate_reg_0[5414]),.o(intermediate_reg_1[2707])); 
mux_module mux_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5413]),.i2(intermediate_reg_0[5412]),.o(intermediate_reg_1[2706]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5411]),.i2(intermediate_reg_0[5410]),.o(intermediate_reg_1[2705]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5409]),.i2(intermediate_reg_0[5408]),.o(intermediate_reg_1[2704])); 
mux_module mux_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5407]),.i2(intermediate_reg_0[5406]),.o(intermediate_reg_1[2703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5405]),.i2(intermediate_reg_0[5404]),.o(intermediate_reg_1[2702]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5403]),.i2(intermediate_reg_0[5402]),.o(intermediate_reg_1[2701]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5401]),.i2(intermediate_reg_0[5400]),.o(intermediate_reg_1[2700])); 
xor_module xor_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5399]),.i2(intermediate_reg_0[5398]),.o(intermediate_reg_1[2699])); 
mux_module mux_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5397]),.i2(intermediate_reg_0[5396]),.o(intermediate_reg_1[2698]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5395]),.i2(intermediate_reg_0[5394]),.o(intermediate_reg_1[2697])); 
mux_module mux_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5393]),.i2(intermediate_reg_0[5392]),.o(intermediate_reg_1[2696]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5391]),.i2(intermediate_reg_0[5390]),.o(intermediate_reg_1[2695])); 
mux_module mux_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5389]),.i2(intermediate_reg_0[5388]),.o(intermediate_reg_1[2694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5387]),.i2(intermediate_reg_0[5386]),.o(intermediate_reg_1[2693]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5385]),.i2(intermediate_reg_0[5384]),.o(intermediate_reg_1[2692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5383]),.i2(intermediate_reg_0[5382]),.o(intermediate_reg_1[2691]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5381]),.i2(intermediate_reg_0[5380]),.o(intermediate_reg_1[2690])); 
mux_module mux_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5379]),.i2(intermediate_reg_0[5378]),.o(intermediate_reg_1[2689]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5377]),.i2(intermediate_reg_0[5376]),.o(intermediate_reg_1[2688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5375]),.i2(intermediate_reg_0[5374]),.o(intermediate_reg_1[2687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5373]),.i2(intermediate_reg_0[5372]),.o(intermediate_reg_1[2686]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5371]),.i2(intermediate_reg_0[5370]),.o(intermediate_reg_1[2685]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5369]),.i2(intermediate_reg_0[5368]),.o(intermediate_reg_1[2684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5367]),.i2(intermediate_reg_0[5366]),.o(intermediate_reg_1[2683]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5365]),.i2(intermediate_reg_0[5364]),.o(intermediate_reg_1[2682])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5363]),.i2(intermediate_reg_0[5362]),.o(intermediate_reg_1[2681]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5361]),.i2(intermediate_reg_0[5360]),.o(intermediate_reg_1[2680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5359]),.i2(intermediate_reg_0[5358]),.o(intermediate_reg_1[2679]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5357]),.i2(intermediate_reg_0[5356]),.o(intermediate_reg_1[2678])); 
xor_module xor_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5355]),.i2(intermediate_reg_0[5354]),.o(intermediate_reg_1[2677])); 
xor_module xor_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5353]),.i2(intermediate_reg_0[5352]),.o(intermediate_reg_1[2676])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5351]),.i2(intermediate_reg_0[5350]),.o(intermediate_reg_1[2675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5349]),.i2(intermediate_reg_0[5348]),.o(intermediate_reg_1[2674]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5347]),.i2(intermediate_reg_0[5346]),.o(intermediate_reg_1[2673])); 
mux_module mux_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5345]),.i2(intermediate_reg_0[5344]),.o(intermediate_reg_1[2672]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5343]),.i2(intermediate_reg_0[5342]),.o(intermediate_reg_1[2671])); 
xor_module xor_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5341]),.i2(intermediate_reg_0[5340]),.o(intermediate_reg_1[2670])); 
xor_module xor_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5339]),.i2(intermediate_reg_0[5338]),.o(intermediate_reg_1[2669])); 
xor_module xor_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5337]),.i2(intermediate_reg_0[5336]),.o(intermediate_reg_1[2668])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5335]),.i2(intermediate_reg_0[5334]),.o(intermediate_reg_1[2667]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5333]),.i2(intermediate_reg_0[5332]),.o(intermediate_reg_1[2666])); 
xor_module xor_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5331]),.i2(intermediate_reg_0[5330]),.o(intermediate_reg_1[2665])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5329]),.i2(intermediate_reg_0[5328]),.o(intermediate_reg_1[2664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5327]),.i2(intermediate_reg_0[5326]),.o(intermediate_reg_1[2663]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5325]),.i2(intermediate_reg_0[5324]),.o(intermediate_reg_1[2662])); 
mux_module mux_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5323]),.i2(intermediate_reg_0[5322]),.o(intermediate_reg_1[2661]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5321]),.i2(intermediate_reg_0[5320]),.o(intermediate_reg_1[2660]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5319]),.i2(intermediate_reg_0[5318]),.o(intermediate_reg_1[2659]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5317]),.i2(intermediate_reg_0[5316]),.o(intermediate_reg_1[2658])); 
xor_module xor_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5315]),.i2(intermediate_reg_0[5314]),.o(intermediate_reg_1[2657])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5313]),.i2(intermediate_reg_0[5312]),.o(intermediate_reg_1[2656])); 
xor_module xor_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5311]),.i2(intermediate_reg_0[5310]),.o(intermediate_reg_1[2655])); 
mux_module mux_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5309]),.i2(intermediate_reg_0[5308]),.o(intermediate_reg_1[2654]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5307]),.i2(intermediate_reg_0[5306]),.o(intermediate_reg_1[2653]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5305]),.i2(intermediate_reg_0[5304]),.o(intermediate_reg_1[2652])); 
mux_module mux_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5303]),.i2(intermediate_reg_0[5302]),.o(intermediate_reg_1[2651]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5301]),.i2(intermediate_reg_0[5300]),.o(intermediate_reg_1[2650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5299]),.i2(intermediate_reg_0[5298]),.o(intermediate_reg_1[2649]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5297]),.i2(intermediate_reg_0[5296]),.o(intermediate_reg_1[2648]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5295]),.i2(intermediate_reg_0[5294]),.o(intermediate_reg_1[2647]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5293]),.i2(intermediate_reg_0[5292]),.o(intermediate_reg_1[2646]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5291]),.i2(intermediate_reg_0[5290]),.o(intermediate_reg_1[2645]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5289]),.i2(intermediate_reg_0[5288]),.o(intermediate_reg_1[2644]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5287]),.i2(intermediate_reg_0[5286]),.o(intermediate_reg_1[2643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5285]),.i2(intermediate_reg_0[5284]),.o(intermediate_reg_1[2642]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5283]),.i2(intermediate_reg_0[5282]),.o(intermediate_reg_1[2641])); 
xor_module xor_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5281]),.i2(intermediate_reg_0[5280]),.o(intermediate_reg_1[2640])); 
mux_module mux_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5279]),.i2(intermediate_reg_0[5278]),.o(intermediate_reg_1[2639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5277]),.i2(intermediate_reg_0[5276]),.o(intermediate_reg_1[2638]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5275]),.i2(intermediate_reg_0[5274]),.o(intermediate_reg_1[2637]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5273]),.i2(intermediate_reg_0[5272]),.o(intermediate_reg_1[2636])); 
mux_module mux_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5271]),.i2(intermediate_reg_0[5270]),.o(intermediate_reg_1[2635]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5269]),.i2(intermediate_reg_0[5268]),.o(intermediate_reg_1[2634])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5267]),.i2(intermediate_reg_0[5266]),.o(intermediate_reg_1[2633]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5265]),.i2(intermediate_reg_0[5264]),.o(intermediate_reg_1[2632])); 
xor_module xor_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5263]),.i2(intermediate_reg_0[5262]),.o(intermediate_reg_1[2631])); 
xor_module xor_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5261]),.i2(intermediate_reg_0[5260]),.o(intermediate_reg_1[2630])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5259]),.i2(intermediate_reg_0[5258]),.o(intermediate_reg_1[2629]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5257]),.i2(intermediate_reg_0[5256]),.o(intermediate_reg_1[2628])); 
xor_module xor_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5255]),.i2(intermediate_reg_0[5254]),.o(intermediate_reg_1[2627])); 
xor_module xor_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5253]),.i2(intermediate_reg_0[5252]),.o(intermediate_reg_1[2626])); 
xor_module xor_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5251]),.i2(intermediate_reg_0[5250]),.o(intermediate_reg_1[2625])); 
mux_module mux_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5249]),.i2(intermediate_reg_0[5248]),.o(intermediate_reg_1[2624]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5247]),.i2(intermediate_reg_0[5246]),.o(intermediate_reg_1[2623])); 
xor_module xor_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5245]),.i2(intermediate_reg_0[5244]),.o(intermediate_reg_1[2622])); 
mux_module mux_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5243]),.i2(intermediate_reg_0[5242]),.o(intermediate_reg_1[2621]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5241]),.i2(intermediate_reg_0[5240]),.o(intermediate_reg_1[2620])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5239]),.i2(intermediate_reg_0[5238]),.o(intermediate_reg_1[2619])); 
mux_module mux_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5237]),.i2(intermediate_reg_0[5236]),.o(intermediate_reg_1[2618]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5235]),.i2(intermediate_reg_0[5234]),.o(intermediate_reg_1[2617]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5233]),.i2(intermediate_reg_0[5232]),.o(intermediate_reg_1[2616]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5231]),.i2(intermediate_reg_0[5230]),.o(intermediate_reg_1[2615])); 
mux_module mux_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5229]),.i2(intermediate_reg_0[5228]),.o(intermediate_reg_1[2614]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5227]),.i2(intermediate_reg_0[5226]),.o(intermediate_reg_1[2613])); 
xor_module xor_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5225]),.i2(intermediate_reg_0[5224]),.o(intermediate_reg_1[2612])); 
xor_module xor_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5223]),.i2(intermediate_reg_0[5222]),.o(intermediate_reg_1[2611])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5221]),.i2(intermediate_reg_0[5220]),.o(intermediate_reg_1[2610])); 
mux_module mux_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5219]),.i2(intermediate_reg_0[5218]),.o(intermediate_reg_1[2609]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5217]),.i2(intermediate_reg_0[5216]),.o(intermediate_reg_1[2608])); 
mux_module mux_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5215]),.i2(intermediate_reg_0[5214]),.o(intermediate_reg_1[2607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5213]),.i2(intermediate_reg_0[5212]),.o(intermediate_reg_1[2606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5211]),.i2(intermediate_reg_0[5210]),.o(intermediate_reg_1[2605]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5209]),.i2(intermediate_reg_0[5208]),.o(intermediate_reg_1[2604])); 
xor_module xor_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5207]),.i2(intermediate_reg_0[5206]),.o(intermediate_reg_1[2603])); 
xor_module xor_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5205]),.i2(intermediate_reg_0[5204]),.o(intermediate_reg_1[2602])); 
xor_module xor_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5203]),.i2(intermediate_reg_0[5202]),.o(intermediate_reg_1[2601])); 
mux_module mux_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5201]),.i2(intermediate_reg_0[5200]),.o(intermediate_reg_1[2600]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5199]),.i2(intermediate_reg_0[5198]),.o(intermediate_reg_1[2599])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5197]),.i2(intermediate_reg_0[5196]),.o(intermediate_reg_1[2598]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5195]),.i2(intermediate_reg_0[5194]),.o(intermediate_reg_1[2597])); 
xor_module xor_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5193]),.i2(intermediate_reg_0[5192]),.o(intermediate_reg_1[2596])); 
xor_module xor_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5191]),.i2(intermediate_reg_0[5190]),.o(intermediate_reg_1[2595])); 
mux_module mux_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5189]),.i2(intermediate_reg_0[5188]),.o(intermediate_reg_1[2594]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5187]),.i2(intermediate_reg_0[5186]),.o(intermediate_reg_1[2593]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5185]),.i2(intermediate_reg_0[5184]),.o(intermediate_reg_1[2592])); 
xor_module xor_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5183]),.i2(intermediate_reg_0[5182]),.o(intermediate_reg_1[2591])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5181]),.i2(intermediate_reg_0[5180]),.o(intermediate_reg_1[2590]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5179]),.i2(intermediate_reg_0[5178]),.o(intermediate_reg_1[2589]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5177]),.i2(intermediate_reg_0[5176]),.o(intermediate_reg_1[2588]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5175]),.i2(intermediate_reg_0[5174]),.o(intermediate_reg_1[2587]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5173]),.i2(intermediate_reg_0[5172]),.o(intermediate_reg_1[2586])); 
xor_module xor_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5171]),.i2(intermediate_reg_0[5170]),.o(intermediate_reg_1[2585])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5169]),.i2(intermediate_reg_0[5168]),.o(intermediate_reg_1[2584])); 
xor_module xor_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5167]),.i2(intermediate_reg_0[5166]),.o(intermediate_reg_1[2583])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5165]),.i2(intermediate_reg_0[5164]),.o(intermediate_reg_1[2582])); 
xor_module xor_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5163]),.i2(intermediate_reg_0[5162]),.o(intermediate_reg_1[2581])); 
mux_module mux_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5161]),.i2(intermediate_reg_0[5160]),.o(intermediate_reg_1[2580]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5159]),.i2(intermediate_reg_0[5158]),.o(intermediate_reg_1[2579]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5157]),.i2(intermediate_reg_0[5156]),.o(intermediate_reg_1[2578])); 
xor_module xor_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5155]),.i2(intermediate_reg_0[5154]),.o(intermediate_reg_1[2577])); 
xor_module xor_module_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5153]),.i2(intermediate_reg_0[5152]),.o(intermediate_reg_1[2576])); 
mux_module mux_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5151]),.i2(intermediate_reg_0[5150]),.o(intermediate_reg_1[2575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5149]),.i2(intermediate_reg_0[5148]),.o(intermediate_reg_1[2574]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5147]),.i2(intermediate_reg_0[5146]),.o(intermediate_reg_1[2573])); 
mux_module mux_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5145]),.i2(intermediate_reg_0[5144]),.o(intermediate_reg_1[2572]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5143]),.i2(intermediate_reg_0[5142]),.o(intermediate_reg_1[2571]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5141]),.i2(intermediate_reg_0[5140]),.o(intermediate_reg_1[2570])); 
mux_module mux_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5139]),.i2(intermediate_reg_0[5138]),.o(intermediate_reg_1[2569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5137]),.i2(intermediate_reg_0[5136]),.o(intermediate_reg_1[2568]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5135]),.i2(intermediate_reg_0[5134]),.o(intermediate_reg_1[2567])); 
xor_module xor_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5133]),.i2(intermediate_reg_0[5132]),.o(intermediate_reg_1[2566])); 
mux_module mux_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5131]),.i2(intermediate_reg_0[5130]),.o(intermediate_reg_1[2565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5129]),.i2(intermediate_reg_0[5128]),.o(intermediate_reg_1[2564]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5127]),.i2(intermediate_reg_0[5126]),.o(intermediate_reg_1[2563]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5125]),.i2(intermediate_reg_0[5124]),.o(intermediate_reg_1[2562]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5123]),.i2(intermediate_reg_0[5122]),.o(intermediate_reg_1[2561])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5121]),.i2(intermediate_reg_0[5120]),.o(intermediate_reg_1[2560]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5119]),.i2(intermediate_reg_0[5118]),.o(intermediate_reg_1[2559])); 
mux_module mux_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5117]),.i2(intermediate_reg_0[5116]),.o(intermediate_reg_1[2558]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5115]),.i2(intermediate_reg_0[5114]),.o(intermediate_reg_1[2557]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5113]),.i2(intermediate_reg_0[5112]),.o(intermediate_reg_1[2556])); 
mux_module mux_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5111]),.i2(intermediate_reg_0[5110]),.o(intermediate_reg_1[2555]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5109]),.i2(intermediate_reg_0[5108]),.o(intermediate_reg_1[2554]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5107]),.i2(intermediate_reg_0[5106]),.o(intermediate_reg_1[2553])); 
xor_module xor_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5105]),.i2(intermediate_reg_0[5104]),.o(intermediate_reg_1[2552])); 
mux_module mux_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5103]),.i2(intermediate_reg_0[5102]),.o(intermediate_reg_1[2551]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5101]),.i2(intermediate_reg_0[5100]),.o(intermediate_reg_1[2550])); 
xor_module xor_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5099]),.i2(intermediate_reg_0[5098]),.o(intermediate_reg_1[2549])); 
xor_module xor_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5097]),.i2(intermediate_reg_0[5096]),.o(intermediate_reg_1[2548])); 
mux_module mux_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5095]),.i2(intermediate_reg_0[5094]),.o(intermediate_reg_1[2547]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5093]),.i2(intermediate_reg_0[5092]),.o(intermediate_reg_1[2546])); 
mux_module mux_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5091]),.i2(intermediate_reg_0[5090]),.o(intermediate_reg_1[2545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5089]),.i2(intermediate_reg_0[5088]),.o(intermediate_reg_1[2544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5087]),.i2(intermediate_reg_0[5086]),.o(intermediate_reg_1[2543]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5085]),.i2(intermediate_reg_0[5084]),.o(intermediate_reg_1[2542]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5083]),.i2(intermediate_reg_0[5082]),.o(intermediate_reg_1[2541])); 
xor_module xor_module_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5081]),.i2(intermediate_reg_0[5080]),.o(intermediate_reg_1[2540])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5079]),.i2(intermediate_reg_0[5078]),.o(intermediate_reg_1[2539]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5077]),.i2(intermediate_reg_0[5076]),.o(intermediate_reg_1[2538])); 
mux_module mux_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5075]),.i2(intermediate_reg_0[5074]),.o(intermediate_reg_1[2537]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5073]),.i2(intermediate_reg_0[5072]),.o(intermediate_reg_1[2536]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5071]),.i2(intermediate_reg_0[5070]),.o(intermediate_reg_1[2535]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5069]),.i2(intermediate_reg_0[5068]),.o(intermediate_reg_1[2534]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5067]),.i2(intermediate_reg_0[5066]),.o(intermediate_reg_1[2533])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5065]),.i2(intermediate_reg_0[5064]),.o(intermediate_reg_1[2532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5063]),.i2(intermediate_reg_0[5062]),.o(intermediate_reg_1[2531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5061]),.i2(intermediate_reg_0[5060]),.o(intermediate_reg_1[2530]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5059]),.i2(intermediate_reg_0[5058]),.o(intermediate_reg_1[2529]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5057]),.i2(intermediate_reg_0[5056]),.o(intermediate_reg_1[2528])); 
mux_module mux_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5055]),.i2(intermediate_reg_0[5054]),.o(intermediate_reg_1[2527]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5053]),.i2(intermediate_reg_0[5052]),.o(intermediate_reg_1[2526]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5051]),.i2(intermediate_reg_0[5050]),.o(intermediate_reg_1[2525])); 
mux_module mux_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5049]),.i2(intermediate_reg_0[5048]),.o(intermediate_reg_1[2524]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5047]),.i2(intermediate_reg_0[5046]),.o(intermediate_reg_1[2523])); 
mux_module mux_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5045]),.i2(intermediate_reg_0[5044]),.o(intermediate_reg_1[2522]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5043]),.i2(intermediate_reg_0[5042]),.o(intermediate_reg_1[2521])); 
mux_module mux_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5041]),.i2(intermediate_reg_0[5040]),.o(intermediate_reg_1[2520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5039]),.i2(intermediate_reg_0[5038]),.o(intermediate_reg_1[2519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5037]),.i2(intermediate_reg_0[5036]),.o(intermediate_reg_1[2518]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5035]),.i2(intermediate_reg_0[5034]),.o(intermediate_reg_1[2517])); 
xor_module xor_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5033]),.i2(intermediate_reg_0[5032]),.o(intermediate_reg_1[2516])); 
xor_module xor_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5031]),.i2(intermediate_reg_0[5030]),.o(intermediate_reg_1[2515])); 
xor_module xor_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5029]),.i2(intermediate_reg_0[5028]),.o(intermediate_reg_1[2514])); 
mux_module mux_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5027]),.i2(intermediate_reg_0[5026]),.o(intermediate_reg_1[2513]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5025]),.i2(intermediate_reg_0[5024]),.o(intermediate_reg_1[2512])); 
xor_module xor_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5023]),.i2(intermediate_reg_0[5022]),.o(intermediate_reg_1[2511])); 
mux_module mux_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5021]),.i2(intermediate_reg_0[5020]),.o(intermediate_reg_1[2510]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5019]),.i2(intermediate_reg_0[5018]),.o(intermediate_reg_1[2509])); 
mux_module mux_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5017]),.i2(intermediate_reg_0[5016]),.o(intermediate_reg_1[2508]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5015]),.i2(intermediate_reg_0[5014]),.o(intermediate_reg_1[2507])); 
xor_module xor_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5013]),.i2(intermediate_reg_0[5012]),.o(intermediate_reg_1[2506])); 
mux_module mux_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5011]),.i2(intermediate_reg_0[5010]),.o(intermediate_reg_1[2505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5009]),.i2(intermediate_reg_0[5008]),.o(intermediate_reg_1[2504]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5007]),.i2(intermediate_reg_0[5006]),.o(intermediate_reg_1[2503]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5005]),.i2(intermediate_reg_0[5004]),.o(intermediate_reg_1[2502])); 
mux_module mux_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5003]),.i2(intermediate_reg_0[5002]),.o(intermediate_reg_1[2501]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5001]),.i2(intermediate_reg_0[5000]),.o(intermediate_reg_1[2500])); 
mux_module mux_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4999]),.i2(intermediate_reg_0[4998]),.o(intermediate_reg_1[2499]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4997]),.i2(intermediate_reg_0[4996]),.o(intermediate_reg_1[2498]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4995]),.i2(intermediate_reg_0[4994]),.o(intermediate_reg_1[2497])); 
xor_module xor_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4993]),.i2(intermediate_reg_0[4992]),.o(intermediate_reg_1[2496])); 
mux_module mux_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4991]),.i2(intermediate_reg_0[4990]),.o(intermediate_reg_1[2495]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4989]),.i2(intermediate_reg_0[4988]),.o(intermediate_reg_1[2494])); 
mux_module mux_module_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4987]),.i2(intermediate_reg_0[4986]),.o(intermediate_reg_1[2493]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4985]),.i2(intermediate_reg_0[4984]),.o(intermediate_reg_1[2492])); 
mux_module mux_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4983]),.i2(intermediate_reg_0[4982]),.o(intermediate_reg_1[2491]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4981]),.i2(intermediate_reg_0[4980]),.o(intermediate_reg_1[2490])); 
xor_module xor_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4979]),.i2(intermediate_reg_0[4978]),.o(intermediate_reg_1[2489])); 
mux_module mux_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4977]),.i2(intermediate_reg_0[4976]),.o(intermediate_reg_1[2488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4975]),.i2(intermediate_reg_0[4974]),.o(intermediate_reg_1[2487]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4973]),.i2(intermediate_reg_0[4972]),.o(intermediate_reg_1[2486])); 
mux_module mux_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4971]),.i2(intermediate_reg_0[4970]),.o(intermediate_reg_1[2485]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4969]),.i2(intermediate_reg_0[4968]),.o(intermediate_reg_1[2484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4967]),.i2(intermediate_reg_0[4966]),.o(intermediate_reg_1[2483]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4965]),.i2(intermediate_reg_0[4964]),.o(intermediate_reg_1[2482])); 
mux_module mux_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4963]),.i2(intermediate_reg_0[4962]),.o(intermediate_reg_1[2481]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4961]),.i2(intermediate_reg_0[4960]),.o(intermediate_reg_1[2480])); 
xor_module xor_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4959]),.i2(intermediate_reg_0[4958]),.o(intermediate_reg_1[2479])); 
xor_module xor_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4957]),.i2(intermediate_reg_0[4956]),.o(intermediate_reg_1[2478])); 
mux_module mux_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4955]),.i2(intermediate_reg_0[4954]),.o(intermediate_reg_1[2477]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4953]),.i2(intermediate_reg_0[4952]),.o(intermediate_reg_1[2476]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4951]),.i2(intermediate_reg_0[4950]),.o(intermediate_reg_1[2475]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4949]),.i2(intermediate_reg_0[4948]),.o(intermediate_reg_1[2474])); 
mux_module mux_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4947]),.i2(intermediate_reg_0[4946]),.o(intermediate_reg_1[2473]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4945]),.i2(intermediate_reg_0[4944]),.o(intermediate_reg_1[2472]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4943]),.i2(intermediate_reg_0[4942]),.o(intermediate_reg_1[2471]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4941]),.i2(intermediate_reg_0[4940]),.o(intermediate_reg_1[2470]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4939]),.i2(intermediate_reg_0[4938]),.o(intermediate_reg_1[2469])); 
xor_module xor_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4937]),.i2(intermediate_reg_0[4936]),.o(intermediate_reg_1[2468])); 
xor_module xor_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4935]),.i2(intermediate_reg_0[4934]),.o(intermediate_reg_1[2467])); 
xor_module xor_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4933]),.i2(intermediate_reg_0[4932]),.o(intermediate_reg_1[2466])); 
xor_module xor_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4931]),.i2(intermediate_reg_0[4930]),.o(intermediate_reg_1[2465])); 
mux_module mux_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4929]),.i2(intermediate_reg_0[4928]),.o(intermediate_reg_1[2464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4927]),.i2(intermediate_reg_0[4926]),.o(intermediate_reg_1[2463]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4925]),.i2(intermediate_reg_0[4924]),.o(intermediate_reg_1[2462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4923]),.i2(intermediate_reg_0[4922]),.o(intermediate_reg_1[2461]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4921]),.i2(intermediate_reg_0[4920]),.o(intermediate_reg_1[2460])); 
xor_module xor_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4919]),.i2(intermediate_reg_0[4918]),.o(intermediate_reg_1[2459])); 
mux_module mux_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4917]),.i2(intermediate_reg_0[4916]),.o(intermediate_reg_1[2458]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4915]),.i2(intermediate_reg_0[4914]),.o(intermediate_reg_1[2457])); 
xor_module xor_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4913]),.i2(intermediate_reg_0[4912]),.o(intermediate_reg_1[2456])); 
xor_module xor_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4911]),.i2(intermediate_reg_0[4910]),.o(intermediate_reg_1[2455])); 
mux_module mux_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4909]),.i2(intermediate_reg_0[4908]),.o(intermediate_reg_1[2454]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4907]),.i2(intermediate_reg_0[4906]),.o(intermediate_reg_1[2453])); 
xor_module xor_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4905]),.i2(intermediate_reg_0[4904]),.o(intermediate_reg_1[2452])); 
xor_module xor_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4903]),.i2(intermediate_reg_0[4902]),.o(intermediate_reg_1[2451])); 
mux_module mux_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4901]),.i2(intermediate_reg_0[4900]),.o(intermediate_reg_1[2450]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4899]),.i2(intermediate_reg_0[4898]),.o(intermediate_reg_1[2449])); 
mux_module mux_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4897]),.i2(intermediate_reg_0[4896]),.o(intermediate_reg_1[2448]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4895]),.i2(intermediate_reg_0[4894]),.o(intermediate_reg_1[2447]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4893]),.i2(intermediate_reg_0[4892]),.o(intermediate_reg_1[2446]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4891]),.i2(intermediate_reg_0[4890]),.o(intermediate_reg_1[2445]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4889]),.i2(intermediate_reg_0[4888]),.o(intermediate_reg_1[2444])); 
xor_module xor_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4887]),.i2(intermediate_reg_0[4886]),.o(intermediate_reg_1[2443])); 
xor_module xor_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4885]),.i2(intermediate_reg_0[4884]),.o(intermediate_reg_1[2442])); 
xor_module xor_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4883]),.i2(intermediate_reg_0[4882]),.o(intermediate_reg_1[2441])); 
xor_module xor_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4881]),.i2(intermediate_reg_0[4880]),.o(intermediate_reg_1[2440])); 
mux_module mux_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4879]),.i2(intermediate_reg_0[4878]),.o(intermediate_reg_1[2439]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4877]),.i2(intermediate_reg_0[4876]),.o(intermediate_reg_1[2438])); 
mux_module mux_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4875]),.i2(intermediate_reg_0[4874]),.o(intermediate_reg_1[2437]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4873]),.i2(intermediate_reg_0[4872]),.o(intermediate_reg_1[2436])); 
xor_module xor_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4871]),.i2(intermediate_reg_0[4870]),.o(intermediate_reg_1[2435])); 
mux_module mux_module_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4869]),.i2(intermediate_reg_0[4868]),.o(intermediate_reg_1[2434]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4867]),.i2(intermediate_reg_0[4866]),.o(intermediate_reg_1[2433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4865]),.i2(intermediate_reg_0[4864]),.o(intermediate_reg_1[2432]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4863]),.i2(intermediate_reg_0[4862]),.o(intermediate_reg_1[2431])); 
xor_module xor_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4861]),.i2(intermediate_reg_0[4860]),.o(intermediate_reg_1[2430])); 
xor_module xor_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4859]),.i2(intermediate_reg_0[4858]),.o(intermediate_reg_1[2429])); 
mux_module mux_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4857]),.i2(intermediate_reg_0[4856]),.o(intermediate_reg_1[2428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4855]),.i2(intermediate_reg_0[4854]),.o(intermediate_reg_1[2427]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4853]),.i2(intermediate_reg_0[4852]),.o(intermediate_reg_1[2426])); 
xor_module xor_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4851]),.i2(intermediate_reg_0[4850]),.o(intermediate_reg_1[2425])); 
mux_module mux_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4849]),.i2(intermediate_reg_0[4848]),.o(intermediate_reg_1[2424]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4847]),.i2(intermediate_reg_0[4846]),.o(intermediate_reg_1[2423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4845]),.i2(intermediate_reg_0[4844]),.o(intermediate_reg_1[2422]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4843]),.i2(intermediate_reg_0[4842]),.o(intermediate_reg_1[2421])); 
xor_module xor_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4841]),.i2(intermediate_reg_0[4840]),.o(intermediate_reg_1[2420])); 
mux_module mux_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4839]),.i2(intermediate_reg_0[4838]),.o(intermediate_reg_1[2419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4837]),.i2(intermediate_reg_0[4836]),.o(intermediate_reg_1[2418]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4835]),.i2(intermediate_reg_0[4834]),.o(intermediate_reg_1[2417])); 
mux_module mux_module_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4833]),.i2(intermediate_reg_0[4832]),.o(intermediate_reg_1[2416]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4831]),.i2(intermediate_reg_0[4830]),.o(intermediate_reg_1[2415])); 
xor_module xor_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4829]),.i2(intermediate_reg_0[4828]),.o(intermediate_reg_1[2414])); 
mux_module mux_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4827]),.i2(intermediate_reg_0[4826]),.o(intermediate_reg_1[2413]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4825]),.i2(intermediate_reg_0[4824]),.o(intermediate_reg_1[2412])); 
xor_module xor_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4823]),.i2(intermediate_reg_0[4822]),.o(intermediate_reg_1[2411])); 
xor_module xor_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4821]),.i2(intermediate_reg_0[4820]),.o(intermediate_reg_1[2410])); 
xor_module xor_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4819]),.i2(intermediate_reg_0[4818]),.o(intermediate_reg_1[2409])); 
mux_module mux_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4817]),.i2(intermediate_reg_0[4816]),.o(intermediate_reg_1[2408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4815]),.i2(intermediate_reg_0[4814]),.o(intermediate_reg_1[2407]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4813]),.i2(intermediate_reg_0[4812]),.o(intermediate_reg_1[2406])); 
mux_module mux_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4811]),.i2(intermediate_reg_0[4810]),.o(intermediate_reg_1[2405]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4809]),.i2(intermediate_reg_0[4808]),.o(intermediate_reg_1[2404])); 
mux_module mux_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4807]),.i2(intermediate_reg_0[4806]),.o(intermediate_reg_1[2403]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4805]),.i2(intermediate_reg_0[4804]),.o(intermediate_reg_1[2402])); 
xor_module xor_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4803]),.i2(intermediate_reg_0[4802]),.o(intermediate_reg_1[2401])); 
mux_module mux_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4801]),.i2(intermediate_reg_0[4800]),.o(intermediate_reg_1[2400]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4799]),.i2(intermediate_reg_0[4798]),.o(intermediate_reg_1[2399])); 
mux_module mux_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4797]),.i2(intermediate_reg_0[4796]),.o(intermediate_reg_1[2398]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4795]),.i2(intermediate_reg_0[4794]),.o(intermediate_reg_1[2397]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4793]),.i2(intermediate_reg_0[4792]),.o(intermediate_reg_1[2396])); 
xor_module xor_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4791]),.i2(intermediate_reg_0[4790]),.o(intermediate_reg_1[2395])); 
mux_module mux_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4789]),.i2(intermediate_reg_0[4788]),.o(intermediate_reg_1[2394]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4787]),.i2(intermediate_reg_0[4786]),.o(intermediate_reg_1[2393])); 
mux_module mux_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4785]),.i2(intermediate_reg_0[4784]),.o(intermediate_reg_1[2392]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4783]),.i2(intermediate_reg_0[4782]),.o(intermediate_reg_1[2391]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4781]),.i2(intermediate_reg_0[4780]),.o(intermediate_reg_1[2390]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4779]),.i2(intermediate_reg_0[4778]),.o(intermediate_reg_1[2389]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4777]),.i2(intermediate_reg_0[4776]),.o(intermediate_reg_1[2388])); 
mux_module mux_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4775]),.i2(intermediate_reg_0[4774]),.o(intermediate_reg_1[2387]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4773]),.i2(intermediate_reg_0[4772]),.o(intermediate_reg_1[2386]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4771]),.i2(intermediate_reg_0[4770]),.o(intermediate_reg_1[2385])); 
xor_module xor_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4769]),.i2(intermediate_reg_0[4768]),.o(intermediate_reg_1[2384])); 
xor_module xor_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4767]),.i2(intermediate_reg_0[4766]),.o(intermediate_reg_1[2383])); 
xor_module xor_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4765]),.i2(intermediate_reg_0[4764]),.o(intermediate_reg_1[2382])); 
xor_module xor_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4763]),.i2(intermediate_reg_0[4762]),.o(intermediate_reg_1[2381])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4761]),.i2(intermediate_reg_0[4760]),.o(intermediate_reg_1[2380]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4759]),.i2(intermediate_reg_0[4758]),.o(intermediate_reg_1[2379])); 
xor_module xor_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4757]),.i2(intermediate_reg_0[4756]),.o(intermediate_reg_1[2378])); 
mux_module mux_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4755]),.i2(intermediate_reg_0[4754]),.o(intermediate_reg_1[2377]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4753]),.i2(intermediate_reg_0[4752]),.o(intermediate_reg_1[2376])); 
xor_module xor_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4751]),.i2(intermediate_reg_0[4750]),.o(intermediate_reg_1[2375])); 
mux_module mux_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4749]),.i2(intermediate_reg_0[4748]),.o(intermediate_reg_1[2374]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4747]),.i2(intermediate_reg_0[4746]),.o(intermediate_reg_1[2373])); 
mux_module mux_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4745]),.i2(intermediate_reg_0[4744]),.o(intermediate_reg_1[2372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4743]),.i2(intermediate_reg_0[4742]),.o(intermediate_reg_1[2371]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4741]),.i2(intermediate_reg_0[4740]),.o(intermediate_reg_1[2370])); 
xor_module xor_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4739]),.i2(intermediate_reg_0[4738]),.o(intermediate_reg_1[2369])); 
mux_module mux_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4737]),.i2(intermediate_reg_0[4736]),.o(intermediate_reg_1[2368]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4735]),.i2(intermediate_reg_0[4734]),.o(intermediate_reg_1[2367])); 
xor_module xor_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4733]),.i2(intermediate_reg_0[4732]),.o(intermediate_reg_1[2366])); 
xor_module xor_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4731]),.i2(intermediate_reg_0[4730]),.o(intermediate_reg_1[2365])); 
mux_module mux_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4729]),.i2(intermediate_reg_0[4728]),.o(intermediate_reg_1[2364]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4727]),.i2(intermediate_reg_0[4726]),.o(intermediate_reg_1[2363]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4725]),.i2(intermediate_reg_0[4724]),.o(intermediate_reg_1[2362])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4723]),.i2(intermediate_reg_0[4722]),.o(intermediate_reg_1[2361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4721]),.i2(intermediate_reg_0[4720]),.o(intermediate_reg_1[2360]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4719]),.i2(intermediate_reg_0[4718]),.o(intermediate_reg_1[2359])); 
mux_module mux_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4717]),.i2(intermediate_reg_0[4716]),.o(intermediate_reg_1[2358]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4715]),.i2(intermediate_reg_0[4714]),.o(intermediate_reg_1[2357])); 
xor_module xor_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4713]),.i2(intermediate_reg_0[4712]),.o(intermediate_reg_1[2356])); 
mux_module mux_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4711]),.i2(intermediate_reg_0[4710]),.o(intermediate_reg_1[2355]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4709]),.i2(intermediate_reg_0[4708]),.o(intermediate_reg_1[2354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4707]),.i2(intermediate_reg_0[4706]),.o(intermediate_reg_1[2353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4705]),.i2(intermediate_reg_0[4704]),.o(intermediate_reg_1[2352]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4703]),.i2(intermediate_reg_0[4702]),.o(intermediate_reg_1[2351])); 
xor_module xor_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4701]),.i2(intermediate_reg_0[4700]),.o(intermediate_reg_1[2350])); 
mux_module mux_module_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4699]),.i2(intermediate_reg_0[4698]),.o(intermediate_reg_1[2349]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4697]),.i2(intermediate_reg_0[4696]),.o(intermediate_reg_1[2348])); 
xor_module xor_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4695]),.i2(intermediate_reg_0[4694]),.o(intermediate_reg_1[2347])); 
mux_module mux_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4693]),.i2(intermediate_reg_0[4692]),.o(intermediate_reg_1[2346]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4691]),.i2(intermediate_reg_0[4690]),.o(intermediate_reg_1[2345])); 
xor_module xor_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4689]),.i2(intermediate_reg_0[4688]),.o(intermediate_reg_1[2344])); 
mux_module mux_module_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4687]),.i2(intermediate_reg_0[4686]),.o(intermediate_reg_1[2343]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4685]),.i2(intermediate_reg_0[4684]),.o(intermediate_reg_1[2342]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4683]),.i2(intermediate_reg_0[4682]),.o(intermediate_reg_1[2341])); 
mux_module mux_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4681]),.i2(intermediate_reg_0[4680]),.o(intermediate_reg_1[2340]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4679]),.i2(intermediate_reg_0[4678]),.o(intermediate_reg_1[2339])); 
xor_module xor_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4677]),.i2(intermediate_reg_0[4676]),.o(intermediate_reg_1[2338])); 
xor_module xor_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4675]),.i2(intermediate_reg_0[4674]),.o(intermediate_reg_1[2337])); 
mux_module mux_module_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4673]),.i2(intermediate_reg_0[4672]),.o(intermediate_reg_1[2336]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4671]),.i2(intermediate_reg_0[4670]),.o(intermediate_reg_1[2335])); 
xor_module xor_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4669]),.i2(intermediate_reg_0[4668]),.o(intermediate_reg_1[2334])); 
xor_module xor_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4667]),.i2(intermediate_reg_0[4666]),.o(intermediate_reg_1[2333])); 
mux_module mux_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4665]),.i2(intermediate_reg_0[4664]),.o(intermediate_reg_1[2332]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4663]),.i2(intermediate_reg_0[4662]),.o(intermediate_reg_1[2331])); 
mux_module mux_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4661]),.i2(intermediate_reg_0[4660]),.o(intermediate_reg_1[2330]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4659]),.i2(intermediate_reg_0[4658]),.o(intermediate_reg_1[2329])); 
xor_module xor_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4657]),.i2(intermediate_reg_0[4656]),.o(intermediate_reg_1[2328])); 
mux_module mux_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4655]),.i2(intermediate_reg_0[4654]),.o(intermediate_reg_1[2327]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4653]),.i2(intermediate_reg_0[4652]),.o(intermediate_reg_1[2326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4651]),.i2(intermediate_reg_0[4650]),.o(intermediate_reg_1[2325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4649]),.i2(intermediate_reg_0[4648]),.o(intermediate_reg_1[2324]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4647]),.i2(intermediate_reg_0[4646]),.o(intermediate_reg_1[2323])); 
xor_module xor_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4645]),.i2(intermediate_reg_0[4644]),.o(intermediate_reg_1[2322])); 
mux_module mux_module_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4643]),.i2(intermediate_reg_0[4642]),.o(intermediate_reg_1[2321]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4641]),.i2(intermediate_reg_0[4640]),.o(intermediate_reg_1[2320])); 
mux_module mux_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4639]),.i2(intermediate_reg_0[4638]),.o(intermediate_reg_1[2319]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4637]),.i2(intermediate_reg_0[4636]),.o(intermediate_reg_1[2318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4635]),.i2(intermediate_reg_0[4634]),.o(intermediate_reg_1[2317]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4633]),.i2(intermediate_reg_0[4632]),.o(intermediate_reg_1[2316])); 
xor_module xor_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4631]),.i2(intermediate_reg_0[4630]),.o(intermediate_reg_1[2315])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4629]),.i2(intermediate_reg_0[4628]),.o(intermediate_reg_1[2314]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4627]),.i2(intermediate_reg_0[4626]),.o(intermediate_reg_1[2313])); 
xor_module xor_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4625]),.i2(intermediate_reg_0[4624]),.o(intermediate_reg_1[2312])); 
mux_module mux_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4623]),.i2(intermediate_reg_0[4622]),.o(intermediate_reg_1[2311]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4621]),.i2(intermediate_reg_0[4620]),.o(intermediate_reg_1[2310])); 
xor_module xor_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4619]),.i2(intermediate_reg_0[4618]),.o(intermediate_reg_1[2309])); 
mux_module mux_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4617]),.i2(intermediate_reg_0[4616]),.o(intermediate_reg_1[2308]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4615]),.i2(intermediate_reg_0[4614]),.o(intermediate_reg_1[2307])); 
mux_module mux_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4613]),.i2(intermediate_reg_0[4612]),.o(intermediate_reg_1[2306]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4611]),.i2(intermediate_reg_0[4610]),.o(intermediate_reg_1[2305])); 
xor_module xor_module_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4609]),.i2(intermediate_reg_0[4608]),.o(intermediate_reg_1[2304])); 
mux_module mux_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4607]),.i2(intermediate_reg_0[4606]),.o(intermediate_reg_1[2303]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4605]),.i2(intermediate_reg_0[4604]),.o(intermediate_reg_1[2302])); 
mux_module mux_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4603]),.i2(intermediate_reg_0[4602]),.o(intermediate_reg_1[2301]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4601]),.i2(intermediate_reg_0[4600]),.o(intermediate_reg_1[2300])); 
mux_module mux_module_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4599]),.i2(intermediate_reg_0[4598]),.o(intermediate_reg_1[2299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4597]),.i2(intermediate_reg_0[4596]),.o(intermediate_reg_1[2298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4595]),.i2(intermediate_reg_0[4594]),.o(intermediate_reg_1[2297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4593]),.i2(intermediate_reg_0[4592]),.o(intermediate_reg_1[2296]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4591]),.i2(intermediate_reg_0[4590]),.o(intermediate_reg_1[2295])); 
xor_module xor_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4589]),.i2(intermediate_reg_0[4588]),.o(intermediate_reg_1[2294])); 
xor_module xor_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4587]),.i2(intermediate_reg_0[4586]),.o(intermediate_reg_1[2293])); 
xor_module xor_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4585]),.i2(intermediate_reg_0[4584]),.o(intermediate_reg_1[2292])); 
mux_module mux_module_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4583]),.i2(intermediate_reg_0[4582]),.o(intermediate_reg_1[2291]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4581]),.i2(intermediate_reg_0[4580]),.o(intermediate_reg_1[2290])); 
xor_module xor_module_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4579]),.i2(intermediate_reg_0[4578]),.o(intermediate_reg_1[2289])); 
xor_module xor_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4577]),.i2(intermediate_reg_0[4576]),.o(intermediate_reg_1[2288])); 
mux_module mux_module_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4575]),.i2(intermediate_reg_0[4574]),.o(intermediate_reg_1[2287]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4573]),.i2(intermediate_reg_0[4572]),.o(intermediate_reg_1[2286])); 
mux_module mux_module_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4571]),.i2(intermediate_reg_0[4570]),.o(intermediate_reg_1[2285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4569]),.i2(intermediate_reg_0[4568]),.o(intermediate_reg_1[2284]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4567]),.i2(intermediate_reg_0[4566]),.o(intermediate_reg_1[2283])); 
mux_module mux_module_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4565]),.i2(intermediate_reg_0[4564]),.o(intermediate_reg_1[2282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4563]),.i2(intermediate_reg_0[4562]),.o(intermediate_reg_1[2281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4561]),.i2(intermediate_reg_0[4560]),.o(intermediate_reg_1[2280]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4559]),.i2(intermediate_reg_0[4558]),.o(intermediate_reg_1[2279])); 
xor_module xor_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4557]),.i2(intermediate_reg_0[4556]),.o(intermediate_reg_1[2278])); 
mux_module mux_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4555]),.i2(intermediate_reg_0[4554]),.o(intermediate_reg_1[2277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4553]),.i2(intermediate_reg_0[4552]),.o(intermediate_reg_1[2276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4551]),.i2(intermediate_reg_0[4550]),.o(intermediate_reg_1[2275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4549]),.i2(intermediate_reg_0[4548]),.o(intermediate_reg_1[2274]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4547]),.i2(intermediate_reg_0[4546]),.o(intermediate_reg_1[2273]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4545]),.i2(intermediate_reg_0[4544]),.o(intermediate_reg_1[2272])); 
mux_module mux_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4543]),.i2(intermediate_reg_0[4542]),.o(intermediate_reg_1[2271]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4541]),.i2(intermediate_reg_0[4540]),.o(intermediate_reg_1[2270])); 
mux_module mux_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4539]),.i2(intermediate_reg_0[4538]),.o(intermediate_reg_1[2269]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4537]),.i2(intermediate_reg_0[4536]),.o(intermediate_reg_1[2268]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4535]),.i2(intermediate_reg_0[4534]),.o(intermediate_reg_1[2267]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4533]),.i2(intermediate_reg_0[4532]),.o(intermediate_reg_1[2266])); 
mux_module mux_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4531]),.i2(intermediate_reg_0[4530]),.o(intermediate_reg_1[2265]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4529]),.i2(intermediate_reg_0[4528]),.o(intermediate_reg_1[2264]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4527]),.i2(intermediate_reg_0[4526]),.o(intermediate_reg_1[2263]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4525]),.i2(intermediate_reg_0[4524]),.o(intermediate_reg_1[2262])); 
mux_module mux_module_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4523]),.i2(intermediate_reg_0[4522]),.o(intermediate_reg_1[2261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4521]),.i2(intermediate_reg_0[4520]),.o(intermediate_reg_1[2260]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4519]),.i2(intermediate_reg_0[4518]),.o(intermediate_reg_1[2259])); 
mux_module mux_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4517]),.i2(intermediate_reg_0[4516]),.o(intermediate_reg_1[2258]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4515]),.i2(intermediate_reg_0[4514]),.o(intermediate_reg_1[2257])); 
mux_module mux_module_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4513]),.i2(intermediate_reg_0[4512]),.o(intermediate_reg_1[2256]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4511]),.i2(intermediate_reg_0[4510]),.o(intermediate_reg_1[2255])); 
xor_module xor_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4509]),.i2(intermediate_reg_0[4508]),.o(intermediate_reg_1[2254])); 
mux_module mux_module_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4507]),.i2(intermediate_reg_0[4506]),.o(intermediate_reg_1[2253]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4505]),.i2(intermediate_reg_0[4504]),.o(intermediate_reg_1[2252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4503]),.i2(intermediate_reg_0[4502]),.o(intermediate_reg_1[2251]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4501]),.i2(intermediate_reg_0[4500]),.o(intermediate_reg_1[2250])); 
mux_module mux_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4499]),.i2(intermediate_reg_0[4498]),.o(intermediate_reg_1[2249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4497]),.i2(intermediate_reg_0[4496]),.o(intermediate_reg_1[2248]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4495]),.i2(intermediate_reg_0[4494]),.o(intermediate_reg_1[2247])); 
xor_module xor_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4493]),.i2(intermediate_reg_0[4492]),.o(intermediate_reg_1[2246])); 
xor_module xor_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4491]),.i2(intermediate_reg_0[4490]),.o(intermediate_reg_1[2245])); 
xor_module xor_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4489]),.i2(intermediate_reg_0[4488]),.o(intermediate_reg_1[2244])); 
mux_module mux_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4487]),.i2(intermediate_reg_0[4486]),.o(intermediate_reg_1[2243]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4485]),.i2(intermediate_reg_0[4484]),.o(intermediate_reg_1[2242])); 
mux_module mux_module_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4483]),.i2(intermediate_reg_0[4482]),.o(intermediate_reg_1[2241]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4481]),.i2(intermediate_reg_0[4480]),.o(intermediate_reg_1[2240])); 
mux_module mux_module_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4479]),.i2(intermediate_reg_0[4478]),.o(intermediate_reg_1[2239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4477]),.i2(intermediate_reg_0[4476]),.o(intermediate_reg_1[2238]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4475]),.i2(intermediate_reg_0[4474]),.o(intermediate_reg_1[2237])); 
xor_module xor_module_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4473]),.i2(intermediate_reg_0[4472]),.o(intermediate_reg_1[2236])); 
xor_module xor_module_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4471]),.i2(intermediate_reg_0[4470]),.o(intermediate_reg_1[2235])); 
mux_module mux_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4469]),.i2(intermediate_reg_0[4468]),.o(intermediate_reg_1[2234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4467]),.i2(intermediate_reg_0[4466]),.o(intermediate_reg_1[2233]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4465]),.i2(intermediate_reg_0[4464]),.o(intermediate_reg_1[2232]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4463]),.i2(intermediate_reg_0[4462]),.o(intermediate_reg_1[2231])); 
mux_module mux_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4461]),.i2(intermediate_reg_0[4460]),.o(intermediate_reg_1[2230]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4459]),.i2(intermediate_reg_0[4458]),.o(intermediate_reg_1[2229])); 
mux_module mux_module_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4457]),.i2(intermediate_reg_0[4456]),.o(intermediate_reg_1[2228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4455]),.i2(intermediate_reg_0[4454]),.o(intermediate_reg_1[2227]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4453]),.i2(intermediate_reg_0[4452]),.o(intermediate_reg_1[2226])); 
mux_module mux_module_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4451]),.i2(intermediate_reg_0[4450]),.o(intermediate_reg_1[2225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4449]),.i2(intermediate_reg_0[4448]),.o(intermediate_reg_1[2224])); 
xor_module xor_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4447]),.i2(intermediate_reg_0[4446]),.o(intermediate_reg_1[2223])); 
mux_module mux_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4445]),.i2(intermediate_reg_0[4444]),.o(intermediate_reg_1[2222]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4443]),.i2(intermediate_reg_0[4442]),.o(intermediate_reg_1[2221])); 
xor_module xor_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4441]),.i2(intermediate_reg_0[4440]),.o(intermediate_reg_1[2220])); 
mux_module mux_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4439]),.i2(intermediate_reg_0[4438]),.o(intermediate_reg_1[2219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4437]),.i2(intermediate_reg_0[4436]),.o(intermediate_reg_1[2218]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4435]),.i2(intermediate_reg_0[4434]),.o(intermediate_reg_1[2217]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4433]),.i2(intermediate_reg_0[4432]),.o(intermediate_reg_1[2216])); 
mux_module mux_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4431]),.i2(intermediate_reg_0[4430]),.o(intermediate_reg_1[2215]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4429]),.i2(intermediate_reg_0[4428]),.o(intermediate_reg_1[2214])); 
xor_module xor_module_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4427]),.i2(intermediate_reg_0[4426]),.o(intermediate_reg_1[2213])); 
mux_module mux_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4425]),.i2(intermediate_reg_0[4424]),.o(intermediate_reg_1[2212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4423]),.i2(intermediate_reg_0[4422]),.o(intermediate_reg_1[2211]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4421]),.i2(intermediate_reg_0[4420]),.o(intermediate_reg_1[2210])); 
xor_module xor_module_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4419]),.i2(intermediate_reg_0[4418]),.o(intermediate_reg_1[2209])); 
mux_module mux_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4417]),.i2(intermediate_reg_0[4416]),.o(intermediate_reg_1[2208]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4415]),.i2(intermediate_reg_0[4414]),.o(intermediate_reg_1[2207])); 
mux_module mux_module_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4413]),.i2(intermediate_reg_0[4412]),.o(intermediate_reg_1[2206]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4411]),.i2(intermediate_reg_0[4410]),.o(intermediate_reg_1[2205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4409]),.i2(intermediate_reg_0[4408]),.o(intermediate_reg_1[2204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4407]),.i2(intermediate_reg_0[4406]),.o(intermediate_reg_1[2203]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4405]),.i2(intermediate_reg_0[4404]),.o(intermediate_reg_1[2202])); 
mux_module mux_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4403]),.i2(intermediate_reg_0[4402]),.o(intermediate_reg_1[2201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4401]),.i2(intermediate_reg_0[4400]),.o(intermediate_reg_1[2200]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4399]),.i2(intermediate_reg_0[4398]),.o(intermediate_reg_1[2199]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4397]),.i2(intermediate_reg_0[4396]),.o(intermediate_reg_1[2198]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4395]),.i2(intermediate_reg_0[4394]),.o(intermediate_reg_1[2197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4393]),.i2(intermediate_reg_0[4392]),.o(intermediate_reg_1[2196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4391]),.i2(intermediate_reg_0[4390]),.o(intermediate_reg_1[2195]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4389]),.i2(intermediate_reg_0[4388]),.o(intermediate_reg_1[2194])); 
mux_module mux_module_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4387]),.i2(intermediate_reg_0[4386]),.o(intermediate_reg_1[2193]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4385]),.i2(intermediate_reg_0[4384]),.o(intermediate_reg_1[2192])); 
xor_module xor_module_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4383]),.i2(intermediate_reg_0[4382]),.o(intermediate_reg_1[2191])); 
mux_module mux_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4381]),.i2(intermediate_reg_0[4380]),.o(intermediate_reg_1[2190]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4379]),.i2(intermediate_reg_0[4378]),.o(intermediate_reg_1[2189])); 
xor_module xor_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4377]),.i2(intermediate_reg_0[4376]),.o(intermediate_reg_1[2188])); 
mux_module mux_module_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4375]),.i2(intermediate_reg_0[4374]),.o(intermediate_reg_1[2187]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4373]),.i2(intermediate_reg_0[4372]),.o(intermediate_reg_1[2186])); 
mux_module mux_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4371]),.i2(intermediate_reg_0[4370]),.o(intermediate_reg_1[2185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4369]),.i2(intermediate_reg_0[4368]),.o(intermediate_reg_1[2184]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4367]),.i2(intermediate_reg_0[4366]),.o(intermediate_reg_1[2183])); 
mux_module mux_module_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4365]),.i2(intermediate_reg_0[4364]),.o(intermediate_reg_1[2182]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4363]),.i2(intermediate_reg_0[4362]),.o(intermediate_reg_1[2181]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4361]),.i2(intermediate_reg_0[4360]),.o(intermediate_reg_1[2180])); 
xor_module xor_module_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4359]),.i2(intermediate_reg_0[4358]),.o(intermediate_reg_1[2179])); 
mux_module mux_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4357]),.i2(intermediate_reg_0[4356]),.o(intermediate_reg_1[2178]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4355]),.i2(intermediate_reg_0[4354]),.o(intermediate_reg_1[2177]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4353]),.i2(intermediate_reg_0[4352]),.o(intermediate_reg_1[2176])); 
xor_module xor_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4351]),.i2(intermediate_reg_0[4350]),.o(intermediate_reg_1[2175])); 
mux_module mux_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4349]),.i2(intermediate_reg_0[4348]),.o(intermediate_reg_1[2174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4347]),.i2(intermediate_reg_0[4346]),.o(intermediate_reg_1[2173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4345]),.i2(intermediate_reg_0[4344]),.o(intermediate_reg_1[2172]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4343]),.i2(intermediate_reg_0[4342]),.o(intermediate_reg_1[2171]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4341]),.i2(intermediate_reg_0[4340]),.o(intermediate_reg_1[2170])); 
mux_module mux_module_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4339]),.i2(intermediate_reg_0[4338]),.o(intermediate_reg_1[2169]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4337]),.i2(intermediate_reg_0[4336]),.o(intermediate_reg_1[2168])); 
xor_module xor_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4335]),.i2(intermediate_reg_0[4334]),.o(intermediate_reg_1[2167])); 
xor_module xor_module_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4333]),.i2(intermediate_reg_0[4332]),.o(intermediate_reg_1[2166])); 
mux_module mux_module_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4331]),.i2(intermediate_reg_0[4330]),.o(intermediate_reg_1[2165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4329]),.i2(intermediate_reg_0[4328]),.o(intermediate_reg_1[2164])); 
mux_module mux_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4327]),.i2(intermediate_reg_0[4326]),.o(intermediate_reg_1[2163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4325]),.i2(intermediate_reg_0[4324]),.o(intermediate_reg_1[2162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4323]),.i2(intermediate_reg_0[4322]),.o(intermediate_reg_1[2161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4321]),.i2(intermediate_reg_0[4320]),.o(intermediate_reg_1[2160]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4319]),.i2(intermediate_reg_0[4318]),.o(intermediate_reg_1[2159])); 
xor_module xor_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4317]),.i2(intermediate_reg_0[4316]),.o(intermediate_reg_1[2158])); 
mux_module mux_module_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4315]),.i2(intermediate_reg_0[4314]),.o(intermediate_reg_1[2157]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4313]),.i2(intermediate_reg_0[4312]),.o(intermediate_reg_1[2156])); 
mux_module mux_module_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4311]),.i2(intermediate_reg_0[4310]),.o(intermediate_reg_1[2155]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4309]),.i2(intermediate_reg_0[4308]),.o(intermediate_reg_1[2154]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4307]),.i2(intermediate_reg_0[4306]),.o(intermediate_reg_1[2153])); 
xor_module xor_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4305]),.i2(intermediate_reg_0[4304]),.o(intermediate_reg_1[2152])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4303]),.i2(intermediate_reg_0[4302]),.o(intermediate_reg_1[2151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4301]),.i2(intermediate_reg_0[4300]),.o(intermediate_reg_1[2150]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4299]),.i2(intermediate_reg_0[4298]),.o(intermediate_reg_1[2149]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4297]),.i2(intermediate_reg_0[4296]),.o(intermediate_reg_1[2148])); 
xor_module xor_module_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4295]),.i2(intermediate_reg_0[4294]),.o(intermediate_reg_1[2147])); 
mux_module mux_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4293]),.i2(intermediate_reg_0[4292]),.o(intermediate_reg_1[2146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4291]),.i2(intermediate_reg_0[4290]),.o(intermediate_reg_1[2145]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4289]),.i2(intermediate_reg_0[4288]),.o(intermediate_reg_1[2144]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4287]),.i2(intermediate_reg_0[4286]),.o(intermediate_reg_1[2143])); 
xor_module xor_module_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4285]),.i2(intermediate_reg_0[4284]),.o(intermediate_reg_1[2142])); 
mux_module mux_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4283]),.i2(intermediate_reg_0[4282]),.o(intermediate_reg_1[2141]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4281]),.i2(intermediate_reg_0[4280]),.o(intermediate_reg_1[2140])); 
xor_module xor_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4279]),.i2(intermediate_reg_0[4278]),.o(intermediate_reg_1[2139])); 
xor_module xor_module_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4277]),.i2(intermediate_reg_0[4276]),.o(intermediate_reg_1[2138])); 
mux_module mux_module_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4275]),.i2(intermediate_reg_0[4274]),.o(intermediate_reg_1[2137]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4273]),.i2(intermediate_reg_0[4272]),.o(intermediate_reg_1[2136]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4271]),.i2(intermediate_reg_0[4270]),.o(intermediate_reg_1[2135])); 
xor_module xor_module_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4269]),.i2(intermediate_reg_0[4268]),.o(intermediate_reg_1[2134])); 
mux_module mux_module_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4267]),.i2(intermediate_reg_0[4266]),.o(intermediate_reg_1[2133]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4265]),.i2(intermediate_reg_0[4264]),.o(intermediate_reg_1[2132])); 
mux_module mux_module_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4263]),.i2(intermediate_reg_0[4262]),.o(intermediate_reg_1[2131]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4261]),.i2(intermediate_reg_0[4260]),.o(intermediate_reg_1[2130])); 
mux_module mux_module_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4259]),.i2(intermediate_reg_0[4258]),.o(intermediate_reg_1[2129]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4257]),.i2(intermediate_reg_0[4256]),.o(intermediate_reg_1[2128])); 
mux_module mux_module_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4255]),.i2(intermediate_reg_0[4254]),.o(intermediate_reg_1[2127]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4253]),.i2(intermediate_reg_0[4252]),.o(intermediate_reg_1[2126])); 
xor_module xor_module_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4251]),.i2(intermediate_reg_0[4250]),.o(intermediate_reg_1[2125])); 
mux_module mux_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4249]),.i2(intermediate_reg_0[4248]),.o(intermediate_reg_1[2124]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4247]),.i2(intermediate_reg_0[4246]),.o(intermediate_reg_1[2123])); 
mux_module mux_module_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4245]),.i2(intermediate_reg_0[4244]),.o(intermediate_reg_1[2122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4243]),.i2(intermediate_reg_0[4242]),.o(intermediate_reg_1[2121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4241]),.i2(intermediate_reg_0[4240]),.o(intermediate_reg_1[2120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4239]),.i2(intermediate_reg_0[4238]),.o(intermediate_reg_1[2119]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4237]),.i2(intermediate_reg_0[4236]),.o(intermediate_reg_1[2118])); 
xor_module xor_module_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4235]),.i2(intermediate_reg_0[4234]),.o(intermediate_reg_1[2117])); 
mux_module mux_module_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4233]),.i2(intermediate_reg_0[4232]),.o(intermediate_reg_1[2116]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4231]),.i2(intermediate_reg_0[4230]),.o(intermediate_reg_1[2115]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4229]),.i2(intermediate_reg_0[4228]),.o(intermediate_reg_1[2114])); 
xor_module xor_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4227]),.i2(intermediate_reg_0[4226]),.o(intermediate_reg_1[2113])); 
mux_module mux_module_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4225]),.i2(intermediate_reg_0[4224]),.o(intermediate_reg_1[2112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4223]),.i2(intermediate_reg_0[4222]),.o(intermediate_reg_1[2111]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4221]),.i2(intermediate_reg_0[4220]),.o(intermediate_reg_1[2110])); 
mux_module mux_module_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4219]),.i2(intermediate_reg_0[4218]),.o(intermediate_reg_1[2109]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4217]),.i2(intermediate_reg_0[4216]),.o(intermediate_reg_1[2108])); 
mux_module mux_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4215]),.i2(intermediate_reg_0[4214]),.o(intermediate_reg_1[2107]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4213]),.i2(intermediate_reg_0[4212]),.o(intermediate_reg_1[2106])); 
mux_module mux_module_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4211]),.i2(intermediate_reg_0[4210]),.o(intermediate_reg_1[2105]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4209]),.i2(intermediate_reg_0[4208]),.o(intermediate_reg_1[2104]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4207]),.i2(intermediate_reg_0[4206]),.o(intermediate_reg_1[2103])); 
xor_module xor_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4205]),.i2(intermediate_reg_0[4204]),.o(intermediate_reg_1[2102])); 
xor_module xor_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4203]),.i2(intermediate_reg_0[4202]),.o(intermediate_reg_1[2101])); 
mux_module mux_module_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4201]),.i2(intermediate_reg_0[4200]),.o(intermediate_reg_1[2100]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4199]),.i2(intermediate_reg_0[4198]),.o(intermediate_reg_1[2099])); 
xor_module xor_module_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4197]),.i2(intermediate_reg_0[4196]),.o(intermediate_reg_1[2098])); 
mux_module mux_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4195]),.i2(intermediate_reg_0[4194]),.o(intermediate_reg_1[2097]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4193]),.i2(intermediate_reg_0[4192]),.o(intermediate_reg_1[2096]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4191]),.i2(intermediate_reg_0[4190]),.o(intermediate_reg_1[2095]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4189]),.i2(intermediate_reg_0[4188]),.o(intermediate_reg_1[2094]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4187]),.i2(intermediate_reg_0[4186]),.o(intermediate_reg_1[2093]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4185]),.i2(intermediate_reg_0[4184]),.o(intermediate_reg_1[2092])); 
mux_module mux_module_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4183]),.i2(intermediate_reg_0[4182]),.o(intermediate_reg_1[2091]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4181]),.i2(intermediate_reg_0[4180]),.o(intermediate_reg_1[2090]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4179]),.i2(intermediate_reg_0[4178]),.o(intermediate_reg_1[2089])); 
mux_module mux_module_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4177]),.i2(intermediate_reg_0[4176]),.o(intermediate_reg_1[2088]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4175]),.i2(intermediate_reg_0[4174]),.o(intermediate_reg_1[2087]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4173]),.i2(intermediate_reg_0[4172]),.o(intermediate_reg_1[2086]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4171]),.i2(intermediate_reg_0[4170]),.o(intermediate_reg_1[2085]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4169]),.i2(intermediate_reg_0[4168]),.o(intermediate_reg_1[2084]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4167]),.i2(intermediate_reg_0[4166]),.o(intermediate_reg_1[2083])); 
xor_module xor_module_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4165]),.i2(intermediate_reg_0[4164]),.o(intermediate_reg_1[2082])); 
xor_module xor_module_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4163]),.i2(intermediate_reg_0[4162]),.o(intermediate_reg_1[2081])); 
mux_module mux_module_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4161]),.i2(intermediate_reg_0[4160]),.o(intermediate_reg_1[2080]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4159]),.i2(intermediate_reg_0[4158]),.o(intermediate_reg_1[2079]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4157]),.i2(intermediate_reg_0[4156]),.o(intermediate_reg_1[2078])); 
mux_module mux_module_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4155]),.i2(intermediate_reg_0[4154]),.o(intermediate_reg_1[2077]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4153]),.i2(intermediate_reg_0[4152]),.o(intermediate_reg_1[2076])); 
mux_module mux_module_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4151]),.i2(intermediate_reg_0[4150]),.o(intermediate_reg_1[2075]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4149]),.i2(intermediate_reg_0[4148]),.o(intermediate_reg_1[2074])); 
xor_module xor_module_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4147]),.i2(intermediate_reg_0[4146]),.o(intermediate_reg_1[2073])); 
xor_module xor_module_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4145]),.i2(intermediate_reg_0[4144]),.o(intermediate_reg_1[2072])); 
mux_module mux_module_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4143]),.i2(intermediate_reg_0[4142]),.o(intermediate_reg_1[2071]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4141]),.i2(intermediate_reg_0[4140]),.o(intermediate_reg_1[2070]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4139]),.i2(intermediate_reg_0[4138]),.o(intermediate_reg_1[2069])); 
mux_module mux_module_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4137]),.i2(intermediate_reg_0[4136]),.o(intermediate_reg_1[2068]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4135]),.i2(intermediate_reg_0[4134]),.o(intermediate_reg_1[2067]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4133]),.i2(intermediate_reg_0[4132]),.o(intermediate_reg_1[2066])); 
xor_module xor_module_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4131]),.i2(intermediate_reg_0[4130]),.o(intermediate_reg_1[2065])); 
xor_module xor_module_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4129]),.i2(intermediate_reg_0[4128]),.o(intermediate_reg_1[2064])); 
xor_module xor_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4127]),.i2(intermediate_reg_0[4126]),.o(intermediate_reg_1[2063])); 
xor_module xor_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4125]),.i2(intermediate_reg_0[4124]),.o(intermediate_reg_1[2062])); 
mux_module mux_module_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4123]),.i2(intermediate_reg_0[4122]),.o(intermediate_reg_1[2061]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4121]),.i2(intermediate_reg_0[4120]),.o(intermediate_reg_1[2060]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4119]),.i2(intermediate_reg_0[4118]),.o(intermediate_reg_1[2059]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4117]),.i2(intermediate_reg_0[4116]),.o(intermediate_reg_1[2058]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4115]),.i2(intermediate_reg_0[4114]),.o(intermediate_reg_1[2057]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4113]),.i2(intermediate_reg_0[4112]),.o(intermediate_reg_1[2056]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4111]),.i2(intermediate_reg_0[4110]),.o(intermediate_reg_1[2055])); 
xor_module xor_module_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4109]),.i2(intermediate_reg_0[4108]),.o(intermediate_reg_1[2054])); 
xor_module xor_module_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4107]),.i2(intermediate_reg_0[4106]),.o(intermediate_reg_1[2053])); 
xor_module xor_module_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4105]),.i2(intermediate_reg_0[4104]),.o(intermediate_reg_1[2052])); 
mux_module mux_module_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4103]),.i2(intermediate_reg_0[4102]),.o(intermediate_reg_1[2051]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4101]),.i2(intermediate_reg_0[4100]),.o(intermediate_reg_1[2050]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4099]),.i2(intermediate_reg_0[4098]),.o(intermediate_reg_1[2049]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4097]),.i2(intermediate_reg_0[4096]),.o(intermediate_reg_1[2048])); 
xor_module xor_module_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4095]),.i2(intermediate_reg_0[4094]),.o(intermediate_reg_1[2047])); 
mux_module mux_module_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4093]),.i2(intermediate_reg_0[4092]),.o(intermediate_reg_1[2046]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4091]),.i2(intermediate_reg_0[4090]),.o(intermediate_reg_1[2045]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4089]),.i2(intermediate_reg_0[4088]),.o(intermediate_reg_1[2044])); 
mux_module mux_module_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4087]),.i2(intermediate_reg_0[4086]),.o(intermediate_reg_1[2043]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4085]),.i2(intermediate_reg_0[4084]),.o(intermediate_reg_1[2042])); 
xor_module xor_module_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4083]),.i2(intermediate_reg_0[4082]),.o(intermediate_reg_1[2041])); 
xor_module xor_module_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4081]),.i2(intermediate_reg_0[4080]),.o(intermediate_reg_1[2040])); 
xor_module xor_module_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4079]),.i2(intermediate_reg_0[4078]),.o(intermediate_reg_1[2039])); 
mux_module mux_module_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4077]),.i2(intermediate_reg_0[4076]),.o(intermediate_reg_1[2038]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4075]),.i2(intermediate_reg_0[4074]),.o(intermediate_reg_1[2037]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4073]),.i2(intermediate_reg_0[4072]),.o(intermediate_reg_1[2036]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4071]),.i2(intermediate_reg_0[4070]),.o(intermediate_reg_1[2035])); 
mux_module mux_module_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4069]),.i2(intermediate_reg_0[4068]),.o(intermediate_reg_1[2034]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4067]),.i2(intermediate_reg_0[4066]),.o(intermediate_reg_1[2033]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4065]),.i2(intermediate_reg_0[4064]),.o(intermediate_reg_1[2032])); 
xor_module xor_module_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4063]),.i2(intermediate_reg_0[4062]),.o(intermediate_reg_1[2031])); 
mux_module mux_module_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4061]),.i2(intermediate_reg_0[4060]),.o(intermediate_reg_1[2030]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4059]),.i2(intermediate_reg_0[4058]),.o(intermediate_reg_1[2029]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4057]),.i2(intermediate_reg_0[4056]),.o(intermediate_reg_1[2028]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4055]),.i2(intermediate_reg_0[4054]),.o(intermediate_reg_1[2027])); 
xor_module xor_module_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4053]),.i2(intermediate_reg_0[4052]),.o(intermediate_reg_1[2026])); 
mux_module mux_module_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4051]),.i2(intermediate_reg_0[4050]),.o(intermediate_reg_1[2025]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4049]),.i2(intermediate_reg_0[4048]),.o(intermediate_reg_1[2024])); 
mux_module mux_module_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4047]),.i2(intermediate_reg_0[4046]),.o(intermediate_reg_1[2023]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4045]),.i2(intermediate_reg_0[4044]),.o(intermediate_reg_1[2022]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4043]),.i2(intermediate_reg_0[4042]),.o(intermediate_reg_1[2021])); 
mux_module mux_module_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4041]),.i2(intermediate_reg_0[4040]),.o(intermediate_reg_1[2020]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4039]),.i2(intermediate_reg_0[4038]),.o(intermediate_reg_1[2019])); 
xor_module xor_module_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4037]),.i2(intermediate_reg_0[4036]),.o(intermediate_reg_1[2018])); 
xor_module xor_module_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4035]),.i2(intermediate_reg_0[4034]),.o(intermediate_reg_1[2017])); 
xor_module xor_module_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4033]),.i2(intermediate_reg_0[4032]),.o(intermediate_reg_1[2016])); 
xor_module xor_module_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4031]),.i2(intermediate_reg_0[4030]),.o(intermediate_reg_1[2015])); 
mux_module mux_module_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4029]),.i2(intermediate_reg_0[4028]),.o(intermediate_reg_1[2014]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4027]),.i2(intermediate_reg_0[4026]),.o(intermediate_reg_1[2013])); 
mux_module mux_module_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4025]),.i2(intermediate_reg_0[4024]),.o(intermediate_reg_1[2012]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4023]),.i2(intermediate_reg_0[4022]),.o(intermediate_reg_1[2011])); 
mux_module mux_module_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4021]),.i2(intermediate_reg_0[4020]),.o(intermediate_reg_1[2010]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4019]),.i2(intermediate_reg_0[4018]),.o(intermediate_reg_1[2009])); 
xor_module xor_module_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4017]),.i2(intermediate_reg_0[4016]),.o(intermediate_reg_1[2008])); 
xor_module xor_module_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4015]),.i2(intermediate_reg_0[4014]),.o(intermediate_reg_1[2007])); 
xor_module xor_module_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4013]),.i2(intermediate_reg_0[4012]),.o(intermediate_reg_1[2006])); 
mux_module mux_module_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4011]),.i2(intermediate_reg_0[4010]),.o(intermediate_reg_1[2005]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4009]),.i2(intermediate_reg_0[4008]),.o(intermediate_reg_1[2004]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4007]),.i2(intermediate_reg_0[4006]),.o(intermediate_reg_1[2003])); 
xor_module xor_module_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4005]),.i2(intermediate_reg_0[4004]),.o(intermediate_reg_1[2002])); 
xor_module xor_module_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4003]),.i2(intermediate_reg_0[4002]),.o(intermediate_reg_1[2001])); 
xor_module xor_module_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4001]),.i2(intermediate_reg_0[4000]),.o(intermediate_reg_1[2000])); 
mux_module mux_module_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3999]),.i2(intermediate_reg_0[3998]),.o(intermediate_reg_1[1999]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3997]),.i2(intermediate_reg_0[3996]),.o(intermediate_reg_1[1998]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3995]),.i2(intermediate_reg_0[3994]),.o(intermediate_reg_1[1997])); 
xor_module xor_module_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3993]),.i2(intermediate_reg_0[3992]),.o(intermediate_reg_1[1996])); 
mux_module mux_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3991]),.i2(intermediate_reg_0[3990]),.o(intermediate_reg_1[1995]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3989]),.i2(intermediate_reg_0[3988]),.o(intermediate_reg_1[1994]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3987]),.i2(intermediate_reg_0[3986]),.o(intermediate_reg_1[1993]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3985]),.i2(intermediate_reg_0[3984]),.o(intermediate_reg_1[1992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3983]),.i2(intermediate_reg_0[3982]),.o(intermediate_reg_1[1991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3981]),.i2(intermediate_reg_0[3980]),.o(intermediate_reg_1[1990]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3979]),.i2(intermediate_reg_0[3978]),.o(intermediate_reg_1[1989]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3977]),.i2(intermediate_reg_0[3976]),.o(intermediate_reg_1[1988])); 
mux_module mux_module_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3975]),.i2(intermediate_reg_0[3974]),.o(intermediate_reg_1[1987]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3973]),.i2(intermediate_reg_0[3972]),.o(intermediate_reg_1[1986]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3971]),.i2(intermediate_reg_0[3970]),.o(intermediate_reg_1[1985]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3969]),.i2(intermediate_reg_0[3968]),.o(intermediate_reg_1[1984]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3967]),.i2(intermediate_reg_0[3966]),.o(intermediate_reg_1[1983]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3965]),.i2(intermediate_reg_0[3964]),.o(intermediate_reg_1[1982])); 
mux_module mux_module_inst_1_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3963]),.i2(intermediate_reg_0[3962]),.o(intermediate_reg_1[1981]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3961]),.i2(intermediate_reg_0[3960]),.o(intermediate_reg_1[1980])); 
mux_module mux_module_inst_1_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3959]),.i2(intermediate_reg_0[3958]),.o(intermediate_reg_1[1979]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3957]),.i2(intermediate_reg_0[3956]),.o(intermediate_reg_1[1978]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3955]),.i2(intermediate_reg_0[3954]),.o(intermediate_reg_1[1977]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3953]),.i2(intermediate_reg_0[3952]),.o(intermediate_reg_1[1976])); 
xor_module xor_module_inst_1_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3951]),.i2(intermediate_reg_0[3950]),.o(intermediate_reg_1[1975])); 
mux_module mux_module_inst_1_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3949]),.i2(intermediate_reg_0[3948]),.o(intermediate_reg_1[1974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3947]),.i2(intermediate_reg_0[3946]),.o(intermediate_reg_1[1973]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3945]),.i2(intermediate_reg_0[3944]),.o(intermediate_reg_1[1972])); 
mux_module mux_module_inst_1_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3943]),.i2(intermediate_reg_0[3942]),.o(intermediate_reg_1[1971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3941]),.i2(intermediate_reg_0[3940]),.o(intermediate_reg_1[1970]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3939]),.i2(intermediate_reg_0[3938]),.o(intermediate_reg_1[1969])); 
xor_module xor_module_inst_1_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3937]),.i2(intermediate_reg_0[3936]),.o(intermediate_reg_1[1968])); 
xor_module xor_module_inst_1_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3935]),.i2(intermediate_reg_0[3934]),.o(intermediate_reg_1[1967])); 
mux_module mux_module_inst_1_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3933]),.i2(intermediate_reg_0[3932]),.o(intermediate_reg_1[1966]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3931]),.i2(intermediate_reg_0[3930]),.o(intermediate_reg_1[1965]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3929]),.i2(intermediate_reg_0[3928]),.o(intermediate_reg_1[1964]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3927]),.i2(intermediate_reg_0[3926]),.o(intermediate_reg_1[1963]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3925]),.i2(intermediate_reg_0[3924]),.o(intermediate_reg_1[1962]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3923]),.i2(intermediate_reg_0[3922]),.o(intermediate_reg_1[1961])); 
mux_module mux_module_inst_1_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3921]),.i2(intermediate_reg_0[3920]),.o(intermediate_reg_1[1960]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3919]),.i2(intermediate_reg_0[3918]),.o(intermediate_reg_1[1959]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3917]),.i2(intermediate_reg_0[3916]),.o(intermediate_reg_1[1958]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3915]),.i2(intermediate_reg_0[3914]),.o(intermediate_reg_1[1957])); 
xor_module xor_module_inst_1_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3913]),.i2(intermediate_reg_0[3912]),.o(intermediate_reg_1[1956])); 
mux_module mux_module_inst_1_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3911]),.i2(intermediate_reg_0[3910]),.o(intermediate_reg_1[1955]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3909]),.i2(intermediate_reg_0[3908]),.o(intermediate_reg_1[1954])); 
mux_module mux_module_inst_1_1344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3907]),.i2(intermediate_reg_0[3906]),.o(intermediate_reg_1[1953]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3905]),.i2(intermediate_reg_0[3904]),.o(intermediate_reg_1[1952])); 
xor_module xor_module_inst_1_1346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3903]),.i2(intermediate_reg_0[3902]),.o(intermediate_reg_1[1951])); 
xor_module xor_module_inst_1_1347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3901]),.i2(intermediate_reg_0[3900]),.o(intermediate_reg_1[1950])); 
xor_module xor_module_inst_1_1348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3899]),.i2(intermediate_reg_0[3898]),.o(intermediate_reg_1[1949])); 
xor_module xor_module_inst_1_1349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3897]),.i2(intermediate_reg_0[3896]),.o(intermediate_reg_1[1948])); 
xor_module xor_module_inst_1_1350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3895]),.i2(intermediate_reg_0[3894]),.o(intermediate_reg_1[1947])); 
xor_module xor_module_inst_1_1351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3893]),.i2(intermediate_reg_0[3892]),.o(intermediate_reg_1[1946])); 
xor_module xor_module_inst_1_1352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3891]),.i2(intermediate_reg_0[3890]),.o(intermediate_reg_1[1945])); 
mux_module mux_module_inst_1_1353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3889]),.i2(intermediate_reg_0[3888]),.o(intermediate_reg_1[1944]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3887]),.i2(intermediate_reg_0[3886]),.o(intermediate_reg_1[1943])); 
xor_module xor_module_inst_1_1355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3885]),.i2(intermediate_reg_0[3884]),.o(intermediate_reg_1[1942])); 
mux_module mux_module_inst_1_1356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3883]),.i2(intermediate_reg_0[3882]),.o(intermediate_reg_1[1941]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3881]),.i2(intermediate_reg_0[3880]),.o(intermediate_reg_1[1940])); 
mux_module mux_module_inst_1_1358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3879]),.i2(intermediate_reg_0[3878]),.o(intermediate_reg_1[1939]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3877]),.i2(intermediate_reg_0[3876]),.o(intermediate_reg_1[1938])); 
mux_module mux_module_inst_1_1360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3875]),.i2(intermediate_reg_0[3874]),.o(intermediate_reg_1[1937]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3873]),.i2(intermediate_reg_0[3872]),.o(intermediate_reg_1[1936]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3871]),.i2(intermediate_reg_0[3870]),.o(intermediate_reg_1[1935]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3869]),.i2(intermediate_reg_0[3868]),.o(intermediate_reg_1[1934]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3867]),.i2(intermediate_reg_0[3866]),.o(intermediate_reg_1[1933])); 
xor_module xor_module_inst_1_1365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3865]),.i2(intermediate_reg_0[3864]),.o(intermediate_reg_1[1932])); 
xor_module xor_module_inst_1_1366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3863]),.i2(intermediate_reg_0[3862]),.o(intermediate_reg_1[1931])); 
mux_module mux_module_inst_1_1367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3861]),.i2(intermediate_reg_0[3860]),.o(intermediate_reg_1[1930]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3859]),.i2(intermediate_reg_0[3858]),.o(intermediate_reg_1[1929]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3857]),.i2(intermediate_reg_0[3856]),.o(intermediate_reg_1[1928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3855]),.i2(intermediate_reg_0[3854]),.o(intermediate_reg_1[1927]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3853]),.i2(intermediate_reg_0[3852]),.o(intermediate_reg_1[1926]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3851]),.i2(intermediate_reg_0[3850]),.o(intermediate_reg_1[1925])); 
mux_module mux_module_inst_1_1373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3849]),.i2(intermediate_reg_0[3848]),.o(intermediate_reg_1[1924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3847]),.i2(intermediate_reg_0[3846]),.o(intermediate_reg_1[1923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3845]),.i2(intermediate_reg_0[3844]),.o(intermediate_reg_1[1922]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3843]),.i2(intermediate_reg_0[3842]),.o(intermediate_reg_1[1921]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3841]),.i2(intermediate_reg_0[3840]),.o(intermediate_reg_1[1920])); 
xor_module xor_module_inst_1_1378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3839]),.i2(intermediate_reg_0[3838]),.o(intermediate_reg_1[1919])); 
xor_module xor_module_inst_1_1379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3837]),.i2(intermediate_reg_0[3836]),.o(intermediate_reg_1[1918])); 
xor_module xor_module_inst_1_1380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3835]),.i2(intermediate_reg_0[3834]),.o(intermediate_reg_1[1917])); 
mux_module mux_module_inst_1_1381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3833]),.i2(intermediate_reg_0[3832]),.o(intermediate_reg_1[1916]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3831]),.i2(intermediate_reg_0[3830]),.o(intermediate_reg_1[1915])); 
mux_module mux_module_inst_1_1383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3829]),.i2(intermediate_reg_0[3828]),.o(intermediate_reg_1[1914]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3827]),.i2(intermediate_reg_0[3826]),.o(intermediate_reg_1[1913])); 
xor_module xor_module_inst_1_1385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3825]),.i2(intermediate_reg_0[3824]),.o(intermediate_reg_1[1912])); 
xor_module xor_module_inst_1_1386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3823]),.i2(intermediate_reg_0[3822]),.o(intermediate_reg_1[1911])); 
xor_module xor_module_inst_1_1387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3821]),.i2(intermediate_reg_0[3820]),.o(intermediate_reg_1[1910])); 
xor_module xor_module_inst_1_1388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3819]),.i2(intermediate_reg_0[3818]),.o(intermediate_reg_1[1909])); 
xor_module xor_module_inst_1_1389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3817]),.i2(intermediate_reg_0[3816]),.o(intermediate_reg_1[1908])); 
xor_module xor_module_inst_1_1390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3815]),.i2(intermediate_reg_0[3814]),.o(intermediate_reg_1[1907])); 
mux_module mux_module_inst_1_1391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3813]),.i2(intermediate_reg_0[3812]),.o(intermediate_reg_1[1906]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3811]),.i2(intermediate_reg_0[3810]),.o(intermediate_reg_1[1905])); 
xor_module xor_module_inst_1_1393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3809]),.i2(intermediate_reg_0[3808]),.o(intermediate_reg_1[1904])); 
xor_module xor_module_inst_1_1394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3807]),.i2(intermediate_reg_0[3806]),.o(intermediate_reg_1[1903])); 
xor_module xor_module_inst_1_1395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3805]),.i2(intermediate_reg_0[3804]),.o(intermediate_reg_1[1902])); 
xor_module xor_module_inst_1_1396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3803]),.i2(intermediate_reg_0[3802]),.o(intermediate_reg_1[1901])); 
mux_module mux_module_inst_1_1397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3801]),.i2(intermediate_reg_0[3800]),.o(intermediate_reg_1[1900]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3799]),.i2(intermediate_reg_0[3798]),.o(intermediate_reg_1[1899])); 
xor_module xor_module_inst_1_1399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3797]),.i2(intermediate_reg_0[3796]),.o(intermediate_reg_1[1898])); 
mux_module mux_module_inst_1_1400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3795]),.i2(intermediate_reg_0[3794]),.o(intermediate_reg_1[1897]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3793]),.i2(intermediate_reg_0[3792]),.o(intermediate_reg_1[1896])); 
mux_module mux_module_inst_1_1402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3791]),.i2(intermediate_reg_0[3790]),.o(intermediate_reg_1[1895]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3789]),.i2(intermediate_reg_0[3788]),.o(intermediate_reg_1[1894]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3787]),.i2(intermediate_reg_0[3786]),.o(intermediate_reg_1[1893])); 
mux_module mux_module_inst_1_1405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3785]),.i2(intermediate_reg_0[3784]),.o(intermediate_reg_1[1892]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3783]),.i2(intermediate_reg_0[3782]),.o(intermediate_reg_1[1891])); 
xor_module xor_module_inst_1_1407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3781]),.i2(intermediate_reg_0[3780]),.o(intermediate_reg_1[1890])); 
mux_module mux_module_inst_1_1408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3779]),.i2(intermediate_reg_0[3778]),.o(intermediate_reg_1[1889]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3777]),.i2(intermediate_reg_0[3776]),.o(intermediate_reg_1[1888]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3775]),.i2(intermediate_reg_0[3774]),.o(intermediate_reg_1[1887]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3773]),.i2(intermediate_reg_0[3772]),.o(intermediate_reg_1[1886]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3771]),.i2(intermediate_reg_0[3770]),.o(intermediate_reg_1[1885]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3769]),.i2(intermediate_reg_0[3768]),.o(intermediate_reg_1[1884])); 
mux_module mux_module_inst_1_1414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3767]),.i2(intermediate_reg_0[3766]),.o(intermediate_reg_1[1883]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3765]),.i2(intermediate_reg_0[3764]),.o(intermediate_reg_1[1882]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3763]),.i2(intermediate_reg_0[3762]),.o(intermediate_reg_1[1881]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3761]),.i2(intermediate_reg_0[3760]),.o(intermediate_reg_1[1880]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3759]),.i2(intermediate_reg_0[3758]),.o(intermediate_reg_1[1879]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3757]),.i2(intermediate_reg_0[3756]),.o(intermediate_reg_1[1878])); 
mux_module mux_module_inst_1_1420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3755]),.i2(intermediate_reg_0[3754]),.o(intermediate_reg_1[1877]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3753]),.i2(intermediate_reg_0[3752]),.o(intermediate_reg_1[1876])); 
xor_module xor_module_inst_1_1422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3751]),.i2(intermediate_reg_0[3750]),.o(intermediate_reg_1[1875])); 
xor_module xor_module_inst_1_1423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3749]),.i2(intermediate_reg_0[3748]),.o(intermediate_reg_1[1874])); 
xor_module xor_module_inst_1_1424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3747]),.i2(intermediate_reg_0[3746]),.o(intermediate_reg_1[1873])); 
mux_module mux_module_inst_1_1425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3745]),.i2(intermediate_reg_0[3744]),.o(intermediate_reg_1[1872]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3743]),.i2(intermediate_reg_0[3742]),.o(intermediate_reg_1[1871]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3741]),.i2(intermediate_reg_0[3740]),.o(intermediate_reg_1[1870]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3739]),.i2(intermediate_reg_0[3738]),.o(intermediate_reg_1[1869])); 
xor_module xor_module_inst_1_1429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3737]),.i2(intermediate_reg_0[3736]),.o(intermediate_reg_1[1868])); 
xor_module xor_module_inst_1_1430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3735]),.i2(intermediate_reg_0[3734]),.o(intermediate_reg_1[1867])); 
mux_module mux_module_inst_1_1431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3733]),.i2(intermediate_reg_0[3732]),.o(intermediate_reg_1[1866]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3731]),.i2(intermediate_reg_0[3730]),.o(intermediate_reg_1[1865]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3729]),.i2(intermediate_reg_0[3728]),.o(intermediate_reg_1[1864])); 
xor_module xor_module_inst_1_1434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3727]),.i2(intermediate_reg_0[3726]),.o(intermediate_reg_1[1863])); 
mux_module mux_module_inst_1_1435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3725]),.i2(intermediate_reg_0[3724]),.o(intermediate_reg_1[1862]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3723]),.i2(intermediate_reg_0[3722]),.o(intermediate_reg_1[1861]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3721]),.i2(intermediate_reg_0[3720]),.o(intermediate_reg_1[1860])); 
xor_module xor_module_inst_1_1438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3719]),.i2(intermediate_reg_0[3718]),.o(intermediate_reg_1[1859])); 
mux_module mux_module_inst_1_1439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3717]),.i2(intermediate_reg_0[3716]),.o(intermediate_reg_1[1858]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3715]),.i2(intermediate_reg_0[3714]),.o(intermediate_reg_1[1857])); 
xor_module xor_module_inst_1_1441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3713]),.i2(intermediate_reg_0[3712]),.o(intermediate_reg_1[1856])); 
xor_module xor_module_inst_1_1442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3711]),.i2(intermediate_reg_0[3710]),.o(intermediate_reg_1[1855])); 
mux_module mux_module_inst_1_1443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3709]),.i2(intermediate_reg_0[3708]),.o(intermediate_reg_1[1854]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3707]),.i2(intermediate_reg_0[3706]),.o(intermediate_reg_1[1853]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3705]),.i2(intermediate_reg_0[3704]),.o(intermediate_reg_1[1852]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3703]),.i2(intermediate_reg_0[3702]),.o(intermediate_reg_1[1851])); 
mux_module mux_module_inst_1_1447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3701]),.i2(intermediate_reg_0[3700]),.o(intermediate_reg_1[1850]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3699]),.i2(intermediate_reg_0[3698]),.o(intermediate_reg_1[1849]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3697]),.i2(intermediate_reg_0[3696]),.o(intermediate_reg_1[1848])); 
mux_module mux_module_inst_1_1450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3695]),.i2(intermediate_reg_0[3694]),.o(intermediate_reg_1[1847]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3693]),.i2(intermediate_reg_0[3692]),.o(intermediate_reg_1[1846])); 
xor_module xor_module_inst_1_1452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3691]),.i2(intermediate_reg_0[3690]),.o(intermediate_reg_1[1845])); 
xor_module xor_module_inst_1_1453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3689]),.i2(intermediate_reg_0[3688]),.o(intermediate_reg_1[1844])); 
xor_module xor_module_inst_1_1454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3687]),.i2(intermediate_reg_0[3686]),.o(intermediate_reg_1[1843])); 
xor_module xor_module_inst_1_1455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3685]),.i2(intermediate_reg_0[3684]),.o(intermediate_reg_1[1842])); 
xor_module xor_module_inst_1_1456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3683]),.i2(intermediate_reg_0[3682]),.o(intermediate_reg_1[1841])); 
mux_module mux_module_inst_1_1457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3681]),.i2(intermediate_reg_0[3680]),.o(intermediate_reg_1[1840]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3679]),.i2(intermediate_reg_0[3678]),.o(intermediate_reg_1[1839]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3677]),.i2(intermediate_reg_0[3676]),.o(intermediate_reg_1[1838]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3675]),.i2(intermediate_reg_0[3674]),.o(intermediate_reg_1[1837])); 
xor_module xor_module_inst_1_1461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3673]),.i2(intermediate_reg_0[3672]),.o(intermediate_reg_1[1836])); 
xor_module xor_module_inst_1_1462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3671]),.i2(intermediate_reg_0[3670]),.o(intermediate_reg_1[1835])); 
xor_module xor_module_inst_1_1463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3669]),.i2(intermediate_reg_0[3668]),.o(intermediate_reg_1[1834])); 
xor_module xor_module_inst_1_1464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3667]),.i2(intermediate_reg_0[3666]),.o(intermediate_reg_1[1833])); 
xor_module xor_module_inst_1_1465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3665]),.i2(intermediate_reg_0[3664]),.o(intermediate_reg_1[1832])); 
xor_module xor_module_inst_1_1466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3663]),.i2(intermediate_reg_0[3662]),.o(intermediate_reg_1[1831])); 
xor_module xor_module_inst_1_1467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3661]),.i2(intermediate_reg_0[3660]),.o(intermediate_reg_1[1830])); 
xor_module xor_module_inst_1_1468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3659]),.i2(intermediate_reg_0[3658]),.o(intermediate_reg_1[1829])); 
mux_module mux_module_inst_1_1469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3657]),.i2(intermediate_reg_0[3656]),.o(intermediate_reg_1[1828]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3655]),.i2(intermediate_reg_0[3654]),.o(intermediate_reg_1[1827])); 
mux_module mux_module_inst_1_1471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3653]),.i2(intermediate_reg_0[3652]),.o(intermediate_reg_1[1826]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3651]),.i2(intermediate_reg_0[3650]),.o(intermediate_reg_1[1825])); 
xor_module xor_module_inst_1_1473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3649]),.i2(intermediate_reg_0[3648]),.o(intermediate_reg_1[1824])); 
mux_module mux_module_inst_1_1474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3647]),.i2(intermediate_reg_0[3646]),.o(intermediate_reg_1[1823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3645]),.i2(intermediate_reg_0[3644]),.o(intermediate_reg_1[1822]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3643]),.i2(intermediate_reg_0[3642]),.o(intermediate_reg_1[1821]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3641]),.i2(intermediate_reg_0[3640]),.o(intermediate_reg_1[1820])); 
mux_module mux_module_inst_1_1478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3639]),.i2(intermediate_reg_0[3638]),.o(intermediate_reg_1[1819]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3637]),.i2(intermediate_reg_0[3636]),.o(intermediate_reg_1[1818])); 
mux_module mux_module_inst_1_1480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3635]),.i2(intermediate_reg_0[3634]),.o(intermediate_reg_1[1817]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3633]),.i2(intermediate_reg_0[3632]),.o(intermediate_reg_1[1816])); 
mux_module mux_module_inst_1_1482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3631]),.i2(intermediate_reg_0[3630]),.o(intermediate_reg_1[1815]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3629]),.i2(intermediate_reg_0[3628]),.o(intermediate_reg_1[1814]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3627]),.i2(intermediate_reg_0[3626]),.o(intermediate_reg_1[1813])); 
xor_module xor_module_inst_1_1485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3625]),.i2(intermediate_reg_0[3624]),.o(intermediate_reg_1[1812])); 
mux_module mux_module_inst_1_1486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3623]),.i2(intermediate_reg_0[3622]),.o(intermediate_reg_1[1811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3621]),.i2(intermediate_reg_0[3620]),.o(intermediate_reg_1[1810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3619]),.i2(intermediate_reg_0[3618]),.o(intermediate_reg_1[1809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3617]),.i2(intermediate_reg_0[3616]),.o(intermediate_reg_1[1808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3615]),.i2(intermediate_reg_0[3614]),.o(intermediate_reg_1[1807]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3613]),.i2(intermediate_reg_0[3612]),.o(intermediate_reg_1[1806])); 
mux_module mux_module_inst_1_1492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3611]),.i2(intermediate_reg_0[3610]),.o(intermediate_reg_1[1805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3609]),.i2(intermediate_reg_0[3608]),.o(intermediate_reg_1[1804]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3607]),.i2(intermediate_reg_0[3606]),.o(intermediate_reg_1[1803]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3605]),.i2(intermediate_reg_0[3604]),.o(intermediate_reg_1[1802])); 
xor_module xor_module_inst_1_1496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3603]),.i2(intermediate_reg_0[3602]),.o(intermediate_reg_1[1801])); 
mux_module mux_module_inst_1_1497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3601]),.i2(intermediate_reg_0[3600]),.o(intermediate_reg_1[1800]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3599]),.i2(intermediate_reg_0[3598]),.o(intermediate_reg_1[1799])); 
mux_module mux_module_inst_1_1499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3597]),.i2(intermediate_reg_0[3596]),.o(intermediate_reg_1[1798]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3595]),.i2(intermediate_reg_0[3594]),.o(intermediate_reg_1[1797]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3593]),.i2(intermediate_reg_0[3592]),.o(intermediate_reg_1[1796]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3591]),.i2(intermediate_reg_0[3590]),.o(intermediate_reg_1[1795]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3589]),.i2(intermediate_reg_0[3588]),.o(intermediate_reg_1[1794]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3587]),.i2(intermediate_reg_0[3586]),.o(intermediate_reg_1[1793]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3585]),.i2(intermediate_reg_0[3584]),.o(intermediate_reg_1[1792]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3583]),.i2(intermediate_reg_0[3582]),.o(intermediate_reg_1[1791])); 
mux_module mux_module_inst_1_1507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3581]),.i2(intermediate_reg_0[3580]),.o(intermediate_reg_1[1790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3579]),.i2(intermediate_reg_0[3578]),.o(intermediate_reg_1[1789]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3577]),.i2(intermediate_reg_0[3576]),.o(intermediate_reg_1[1788]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3575]),.i2(intermediate_reg_0[3574]),.o(intermediate_reg_1[1787]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3573]),.i2(intermediate_reg_0[3572]),.o(intermediate_reg_1[1786])); 
mux_module mux_module_inst_1_1512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3571]),.i2(intermediate_reg_0[3570]),.o(intermediate_reg_1[1785]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3569]),.i2(intermediate_reg_0[3568]),.o(intermediate_reg_1[1784]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3567]),.i2(intermediate_reg_0[3566]),.o(intermediate_reg_1[1783])); 
xor_module xor_module_inst_1_1515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3565]),.i2(intermediate_reg_0[3564]),.o(intermediate_reg_1[1782])); 
mux_module mux_module_inst_1_1516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3563]),.i2(intermediate_reg_0[3562]),.o(intermediate_reg_1[1781]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3561]),.i2(intermediate_reg_0[3560]),.o(intermediate_reg_1[1780])); 
xor_module xor_module_inst_1_1518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3559]),.i2(intermediate_reg_0[3558]),.o(intermediate_reg_1[1779])); 
xor_module xor_module_inst_1_1519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3557]),.i2(intermediate_reg_0[3556]),.o(intermediate_reg_1[1778])); 
xor_module xor_module_inst_1_1520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3555]),.i2(intermediate_reg_0[3554]),.o(intermediate_reg_1[1777])); 
xor_module xor_module_inst_1_1521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3553]),.i2(intermediate_reg_0[3552]),.o(intermediate_reg_1[1776])); 
xor_module xor_module_inst_1_1522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3551]),.i2(intermediate_reg_0[3550]),.o(intermediate_reg_1[1775])); 
mux_module mux_module_inst_1_1523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3549]),.i2(intermediate_reg_0[3548]),.o(intermediate_reg_1[1774]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3547]),.i2(intermediate_reg_0[3546]),.o(intermediate_reg_1[1773])); 
mux_module mux_module_inst_1_1525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3545]),.i2(intermediate_reg_0[3544]),.o(intermediate_reg_1[1772]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3543]),.i2(intermediate_reg_0[3542]),.o(intermediate_reg_1[1771])); 
xor_module xor_module_inst_1_1527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3541]),.i2(intermediate_reg_0[3540]),.o(intermediate_reg_1[1770])); 
mux_module mux_module_inst_1_1528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3539]),.i2(intermediate_reg_0[3538]),.o(intermediate_reg_1[1769]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3537]),.i2(intermediate_reg_0[3536]),.o(intermediate_reg_1[1768])); 
mux_module mux_module_inst_1_1530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3535]),.i2(intermediate_reg_0[3534]),.o(intermediate_reg_1[1767]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3533]),.i2(intermediate_reg_0[3532]),.o(intermediate_reg_1[1766])); 
mux_module mux_module_inst_1_1532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3531]),.i2(intermediate_reg_0[3530]),.o(intermediate_reg_1[1765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3529]),.i2(intermediate_reg_0[3528]),.o(intermediate_reg_1[1764]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3527]),.i2(intermediate_reg_0[3526]),.o(intermediate_reg_1[1763])); 
mux_module mux_module_inst_1_1535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3525]),.i2(intermediate_reg_0[3524]),.o(intermediate_reg_1[1762]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3523]),.i2(intermediate_reg_0[3522]),.o(intermediate_reg_1[1761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3521]),.i2(intermediate_reg_0[3520]),.o(intermediate_reg_1[1760]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3519]),.i2(intermediate_reg_0[3518]),.o(intermediate_reg_1[1759])); 
xor_module xor_module_inst_1_1539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3517]),.i2(intermediate_reg_0[3516]),.o(intermediate_reg_1[1758])); 
xor_module xor_module_inst_1_1540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3515]),.i2(intermediate_reg_0[3514]),.o(intermediate_reg_1[1757])); 
xor_module xor_module_inst_1_1541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3513]),.i2(intermediate_reg_0[3512]),.o(intermediate_reg_1[1756])); 
mux_module mux_module_inst_1_1542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3511]),.i2(intermediate_reg_0[3510]),.o(intermediate_reg_1[1755]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3509]),.i2(intermediate_reg_0[3508]),.o(intermediate_reg_1[1754]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3507]),.i2(intermediate_reg_0[3506]),.o(intermediate_reg_1[1753])); 
mux_module mux_module_inst_1_1545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3505]),.i2(intermediate_reg_0[3504]),.o(intermediate_reg_1[1752]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3503]),.i2(intermediate_reg_0[3502]),.o(intermediate_reg_1[1751])); 
mux_module mux_module_inst_1_1547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3501]),.i2(intermediate_reg_0[3500]),.o(intermediate_reg_1[1750]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3499]),.i2(intermediate_reg_0[3498]),.o(intermediate_reg_1[1749]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3497]),.i2(intermediate_reg_0[3496]),.o(intermediate_reg_1[1748]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3495]),.i2(intermediate_reg_0[3494]),.o(intermediate_reg_1[1747]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3493]),.i2(intermediate_reg_0[3492]),.o(intermediate_reg_1[1746])); 
xor_module xor_module_inst_1_1552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3491]),.i2(intermediate_reg_0[3490]),.o(intermediate_reg_1[1745])); 
mux_module mux_module_inst_1_1553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3489]),.i2(intermediate_reg_0[3488]),.o(intermediate_reg_1[1744]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3487]),.i2(intermediate_reg_0[3486]),.o(intermediate_reg_1[1743])); 
xor_module xor_module_inst_1_1555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3485]),.i2(intermediate_reg_0[3484]),.o(intermediate_reg_1[1742])); 
mux_module mux_module_inst_1_1556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3483]),.i2(intermediate_reg_0[3482]),.o(intermediate_reg_1[1741]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3481]),.i2(intermediate_reg_0[3480]),.o(intermediate_reg_1[1740]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3479]),.i2(intermediate_reg_0[3478]),.o(intermediate_reg_1[1739]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3477]),.i2(intermediate_reg_0[3476]),.o(intermediate_reg_1[1738])); 
mux_module mux_module_inst_1_1560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3475]),.i2(intermediate_reg_0[3474]),.o(intermediate_reg_1[1737]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3473]),.i2(intermediate_reg_0[3472]),.o(intermediate_reg_1[1736])); 
xor_module xor_module_inst_1_1562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3471]),.i2(intermediate_reg_0[3470]),.o(intermediate_reg_1[1735])); 
xor_module xor_module_inst_1_1563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3469]),.i2(intermediate_reg_0[3468]),.o(intermediate_reg_1[1734])); 
xor_module xor_module_inst_1_1564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3467]),.i2(intermediate_reg_0[3466]),.o(intermediate_reg_1[1733])); 
xor_module xor_module_inst_1_1565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3465]),.i2(intermediate_reg_0[3464]),.o(intermediate_reg_1[1732])); 
mux_module mux_module_inst_1_1566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3463]),.i2(intermediate_reg_0[3462]),.o(intermediate_reg_1[1731]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3461]),.i2(intermediate_reg_0[3460]),.o(intermediate_reg_1[1730])); 
mux_module mux_module_inst_1_1568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3459]),.i2(intermediate_reg_0[3458]),.o(intermediate_reg_1[1729]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3457]),.i2(intermediate_reg_0[3456]),.o(intermediate_reg_1[1728])); 
xor_module xor_module_inst_1_1570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3455]),.i2(intermediate_reg_0[3454]),.o(intermediate_reg_1[1727])); 
mux_module mux_module_inst_1_1571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3453]),.i2(intermediate_reg_0[3452]),.o(intermediate_reg_1[1726]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3451]),.i2(intermediate_reg_0[3450]),.o(intermediate_reg_1[1725])); 
mux_module mux_module_inst_1_1573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3449]),.i2(intermediate_reg_0[3448]),.o(intermediate_reg_1[1724]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3447]),.i2(intermediate_reg_0[3446]),.o(intermediate_reg_1[1723])); 
xor_module xor_module_inst_1_1575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3445]),.i2(intermediate_reg_0[3444]),.o(intermediate_reg_1[1722])); 
xor_module xor_module_inst_1_1576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3443]),.i2(intermediate_reg_0[3442]),.o(intermediate_reg_1[1721])); 
mux_module mux_module_inst_1_1577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3441]),.i2(intermediate_reg_0[3440]),.o(intermediate_reg_1[1720]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3439]),.i2(intermediate_reg_0[3438]),.o(intermediate_reg_1[1719]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3437]),.i2(intermediate_reg_0[3436]),.o(intermediate_reg_1[1718])); 
xor_module xor_module_inst_1_1580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3435]),.i2(intermediate_reg_0[3434]),.o(intermediate_reg_1[1717])); 
mux_module mux_module_inst_1_1581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3433]),.i2(intermediate_reg_0[3432]),.o(intermediate_reg_1[1716]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3431]),.i2(intermediate_reg_0[3430]),.o(intermediate_reg_1[1715])); 
mux_module mux_module_inst_1_1583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3429]),.i2(intermediate_reg_0[3428]),.o(intermediate_reg_1[1714]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3427]),.i2(intermediate_reg_0[3426]),.o(intermediate_reg_1[1713]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3425]),.i2(intermediate_reg_0[3424]),.o(intermediate_reg_1[1712])); 
xor_module xor_module_inst_1_1586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3423]),.i2(intermediate_reg_0[3422]),.o(intermediate_reg_1[1711])); 
mux_module mux_module_inst_1_1587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3421]),.i2(intermediate_reg_0[3420]),.o(intermediate_reg_1[1710]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3419]),.i2(intermediate_reg_0[3418]),.o(intermediate_reg_1[1709])); 
mux_module mux_module_inst_1_1589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3417]),.i2(intermediate_reg_0[3416]),.o(intermediate_reg_1[1708]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3415]),.i2(intermediate_reg_0[3414]),.o(intermediate_reg_1[1707])); 
xor_module xor_module_inst_1_1591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3413]),.i2(intermediate_reg_0[3412]),.o(intermediate_reg_1[1706])); 
mux_module mux_module_inst_1_1592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3411]),.i2(intermediate_reg_0[3410]),.o(intermediate_reg_1[1705]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3409]),.i2(intermediate_reg_0[3408]),.o(intermediate_reg_1[1704])); 
xor_module xor_module_inst_1_1594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3407]),.i2(intermediate_reg_0[3406]),.o(intermediate_reg_1[1703])); 
xor_module xor_module_inst_1_1595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3405]),.i2(intermediate_reg_0[3404]),.o(intermediate_reg_1[1702])); 
mux_module mux_module_inst_1_1596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3403]),.i2(intermediate_reg_0[3402]),.o(intermediate_reg_1[1701]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3401]),.i2(intermediate_reg_0[3400]),.o(intermediate_reg_1[1700]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3399]),.i2(intermediate_reg_0[3398]),.o(intermediate_reg_1[1699]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3397]),.i2(intermediate_reg_0[3396]),.o(intermediate_reg_1[1698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3395]),.i2(intermediate_reg_0[3394]),.o(intermediate_reg_1[1697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3393]),.i2(intermediate_reg_0[3392]),.o(intermediate_reg_1[1696]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3391]),.i2(intermediate_reg_0[3390]),.o(intermediate_reg_1[1695])); 
mux_module mux_module_inst_1_1603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3389]),.i2(intermediate_reg_0[3388]),.o(intermediate_reg_1[1694]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3387]),.i2(intermediate_reg_0[3386]),.o(intermediate_reg_1[1693])); 
xor_module xor_module_inst_1_1605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3385]),.i2(intermediate_reg_0[3384]),.o(intermediate_reg_1[1692])); 
mux_module mux_module_inst_1_1606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3383]),.i2(intermediate_reg_0[3382]),.o(intermediate_reg_1[1691]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3381]),.i2(intermediate_reg_0[3380]),.o(intermediate_reg_1[1690])); 
xor_module xor_module_inst_1_1608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3379]),.i2(intermediate_reg_0[3378]),.o(intermediate_reg_1[1689])); 
mux_module mux_module_inst_1_1609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3377]),.i2(intermediate_reg_0[3376]),.o(intermediate_reg_1[1688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3375]),.i2(intermediate_reg_0[3374]),.o(intermediate_reg_1[1687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3373]),.i2(intermediate_reg_0[3372]),.o(intermediate_reg_1[1686]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3371]),.i2(intermediate_reg_0[3370]),.o(intermediate_reg_1[1685])); 
xor_module xor_module_inst_1_1613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3369]),.i2(intermediate_reg_0[3368]),.o(intermediate_reg_1[1684])); 
xor_module xor_module_inst_1_1614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3367]),.i2(intermediate_reg_0[3366]),.o(intermediate_reg_1[1683])); 
mux_module mux_module_inst_1_1615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3365]),.i2(intermediate_reg_0[3364]),.o(intermediate_reg_1[1682]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3363]),.i2(intermediate_reg_0[3362]),.o(intermediate_reg_1[1681]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3361]),.i2(intermediate_reg_0[3360]),.o(intermediate_reg_1[1680])); 
mux_module mux_module_inst_1_1618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3359]),.i2(intermediate_reg_0[3358]),.o(intermediate_reg_1[1679]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3357]),.i2(intermediate_reg_0[3356]),.o(intermediate_reg_1[1678])); 
mux_module mux_module_inst_1_1620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3355]),.i2(intermediate_reg_0[3354]),.o(intermediate_reg_1[1677]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3353]),.i2(intermediate_reg_0[3352]),.o(intermediate_reg_1[1676]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3351]),.i2(intermediate_reg_0[3350]),.o(intermediate_reg_1[1675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3349]),.i2(intermediate_reg_0[3348]),.o(intermediate_reg_1[1674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3347]),.i2(intermediate_reg_0[3346]),.o(intermediate_reg_1[1673]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3345]),.i2(intermediate_reg_0[3344]),.o(intermediate_reg_1[1672])); 
xor_module xor_module_inst_1_1626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3343]),.i2(intermediate_reg_0[3342]),.o(intermediate_reg_1[1671])); 
xor_module xor_module_inst_1_1627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3341]),.i2(intermediate_reg_0[3340]),.o(intermediate_reg_1[1670])); 
mux_module mux_module_inst_1_1628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3339]),.i2(intermediate_reg_0[3338]),.o(intermediate_reg_1[1669]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3337]),.i2(intermediate_reg_0[3336]),.o(intermediate_reg_1[1668]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3335]),.i2(intermediate_reg_0[3334]),.o(intermediate_reg_1[1667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3333]),.i2(intermediate_reg_0[3332]),.o(intermediate_reg_1[1666]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3331]),.i2(intermediate_reg_0[3330]),.o(intermediate_reg_1[1665])); 
mux_module mux_module_inst_1_1633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3329]),.i2(intermediate_reg_0[3328]),.o(intermediate_reg_1[1664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3327]),.i2(intermediate_reg_0[3326]),.o(intermediate_reg_1[1663]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3325]),.i2(intermediate_reg_0[3324]),.o(intermediate_reg_1[1662])); 
mux_module mux_module_inst_1_1636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3323]),.i2(intermediate_reg_0[3322]),.o(intermediate_reg_1[1661]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3321]),.i2(intermediate_reg_0[3320]),.o(intermediate_reg_1[1660])); 
mux_module mux_module_inst_1_1638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3319]),.i2(intermediate_reg_0[3318]),.o(intermediate_reg_1[1659]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3317]),.i2(intermediate_reg_0[3316]),.o(intermediate_reg_1[1658])); 
mux_module mux_module_inst_1_1640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3315]),.i2(intermediate_reg_0[3314]),.o(intermediate_reg_1[1657]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3313]),.i2(intermediate_reg_0[3312]),.o(intermediate_reg_1[1656])); 
mux_module mux_module_inst_1_1642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3311]),.i2(intermediate_reg_0[3310]),.o(intermediate_reg_1[1655]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3309]),.i2(intermediate_reg_0[3308]),.o(intermediate_reg_1[1654])); 
xor_module xor_module_inst_1_1644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3307]),.i2(intermediate_reg_0[3306]),.o(intermediate_reg_1[1653])); 
xor_module xor_module_inst_1_1645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3305]),.i2(intermediate_reg_0[3304]),.o(intermediate_reg_1[1652])); 
mux_module mux_module_inst_1_1646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3303]),.i2(intermediate_reg_0[3302]),.o(intermediate_reg_1[1651]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3301]),.i2(intermediate_reg_0[3300]),.o(intermediate_reg_1[1650]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3299]),.i2(intermediate_reg_0[3298]),.o(intermediate_reg_1[1649])); 
xor_module xor_module_inst_1_1649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3297]),.i2(intermediate_reg_0[3296]),.o(intermediate_reg_1[1648])); 
xor_module xor_module_inst_1_1650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3295]),.i2(intermediate_reg_0[3294]),.o(intermediate_reg_1[1647])); 
mux_module mux_module_inst_1_1651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3293]),.i2(intermediate_reg_0[3292]),.o(intermediate_reg_1[1646]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3291]),.i2(intermediate_reg_0[3290]),.o(intermediate_reg_1[1645])); 
xor_module xor_module_inst_1_1653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3289]),.i2(intermediate_reg_0[3288]),.o(intermediate_reg_1[1644])); 
xor_module xor_module_inst_1_1654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3287]),.i2(intermediate_reg_0[3286]),.o(intermediate_reg_1[1643])); 
xor_module xor_module_inst_1_1655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3285]),.i2(intermediate_reg_0[3284]),.o(intermediate_reg_1[1642])); 
xor_module xor_module_inst_1_1656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3283]),.i2(intermediate_reg_0[3282]),.o(intermediate_reg_1[1641])); 
xor_module xor_module_inst_1_1657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3281]),.i2(intermediate_reg_0[3280]),.o(intermediate_reg_1[1640])); 
xor_module xor_module_inst_1_1658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3279]),.i2(intermediate_reg_0[3278]),.o(intermediate_reg_1[1639])); 
xor_module xor_module_inst_1_1659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3277]),.i2(intermediate_reg_0[3276]),.o(intermediate_reg_1[1638])); 
xor_module xor_module_inst_1_1660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3275]),.i2(intermediate_reg_0[3274]),.o(intermediate_reg_1[1637])); 
mux_module mux_module_inst_1_1661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3273]),.i2(intermediate_reg_0[3272]),.o(intermediate_reg_1[1636]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3271]),.i2(intermediate_reg_0[3270]),.o(intermediate_reg_1[1635]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3269]),.i2(intermediate_reg_0[3268]),.o(intermediate_reg_1[1634]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3267]),.i2(intermediate_reg_0[3266]),.o(intermediate_reg_1[1633]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3265]),.i2(intermediate_reg_0[3264]),.o(intermediate_reg_1[1632]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3263]),.i2(intermediate_reg_0[3262]),.o(intermediate_reg_1[1631])); 
mux_module mux_module_inst_1_1667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3261]),.i2(intermediate_reg_0[3260]),.o(intermediate_reg_1[1630]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3259]),.i2(intermediate_reg_0[3258]),.o(intermediate_reg_1[1629]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3257]),.i2(intermediate_reg_0[3256]),.o(intermediate_reg_1[1628]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3255]),.i2(intermediate_reg_0[3254]),.o(intermediate_reg_1[1627]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3253]),.i2(intermediate_reg_0[3252]),.o(intermediate_reg_1[1626]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3251]),.i2(intermediate_reg_0[3250]),.o(intermediate_reg_1[1625]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3249]),.i2(intermediate_reg_0[3248]),.o(intermediate_reg_1[1624]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3247]),.i2(intermediate_reg_0[3246]),.o(intermediate_reg_1[1623]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3245]),.i2(intermediate_reg_0[3244]),.o(intermediate_reg_1[1622])); 
mux_module mux_module_inst_1_1676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3243]),.i2(intermediate_reg_0[3242]),.o(intermediate_reg_1[1621]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3241]),.i2(intermediate_reg_0[3240]),.o(intermediate_reg_1[1620])); 
xor_module xor_module_inst_1_1678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3239]),.i2(intermediate_reg_0[3238]),.o(intermediate_reg_1[1619])); 
mux_module mux_module_inst_1_1679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3237]),.i2(intermediate_reg_0[3236]),.o(intermediate_reg_1[1618]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3235]),.i2(intermediate_reg_0[3234]),.o(intermediate_reg_1[1617])); 
mux_module mux_module_inst_1_1681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3233]),.i2(intermediate_reg_0[3232]),.o(intermediate_reg_1[1616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3231]),.i2(intermediate_reg_0[3230]),.o(intermediate_reg_1[1615]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3229]),.i2(intermediate_reg_0[3228]),.o(intermediate_reg_1[1614])); 
mux_module mux_module_inst_1_1684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3227]),.i2(intermediate_reg_0[3226]),.o(intermediate_reg_1[1613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3225]),.i2(intermediate_reg_0[3224]),.o(intermediate_reg_1[1612]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3223]),.i2(intermediate_reg_0[3222]),.o(intermediate_reg_1[1611]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3221]),.i2(intermediate_reg_0[3220]),.o(intermediate_reg_1[1610]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3219]),.i2(intermediate_reg_0[3218]),.o(intermediate_reg_1[1609])); 
xor_module xor_module_inst_1_1689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3217]),.i2(intermediate_reg_0[3216]),.o(intermediate_reg_1[1608])); 
xor_module xor_module_inst_1_1690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3215]),.i2(intermediate_reg_0[3214]),.o(intermediate_reg_1[1607])); 
mux_module mux_module_inst_1_1691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3213]),.i2(intermediate_reg_0[3212]),.o(intermediate_reg_1[1606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3211]),.i2(intermediate_reg_0[3210]),.o(intermediate_reg_1[1605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3209]),.i2(intermediate_reg_0[3208]),.o(intermediate_reg_1[1604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3207]),.i2(intermediate_reg_0[3206]),.o(intermediate_reg_1[1603]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3205]),.i2(intermediate_reg_0[3204]),.o(intermediate_reg_1[1602])); 
xor_module xor_module_inst_1_1696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3203]),.i2(intermediate_reg_0[3202]),.o(intermediate_reg_1[1601])); 
mux_module mux_module_inst_1_1697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3201]),.i2(intermediate_reg_0[3200]),.o(intermediate_reg_1[1600]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3199]),.i2(intermediate_reg_0[3198]),.o(intermediate_reg_1[1599]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3197]),.i2(intermediate_reg_0[3196]),.o(intermediate_reg_1[1598]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3195]),.i2(intermediate_reg_0[3194]),.o(intermediate_reg_1[1597]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3193]),.i2(intermediate_reg_0[3192]),.o(intermediate_reg_1[1596]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3191]),.i2(intermediate_reg_0[3190]),.o(intermediate_reg_1[1595]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3189]),.i2(intermediate_reg_0[3188]),.o(intermediate_reg_1[1594]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3187]),.i2(intermediate_reg_0[3186]),.o(intermediate_reg_1[1593]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3185]),.i2(intermediate_reg_0[3184]),.o(intermediate_reg_1[1592]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3183]),.i2(intermediate_reg_0[3182]),.o(intermediate_reg_1[1591])); 
mux_module mux_module_inst_1_1707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3181]),.i2(intermediate_reg_0[3180]),.o(intermediate_reg_1[1590]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3179]),.i2(intermediate_reg_0[3178]),.o(intermediate_reg_1[1589])); 
mux_module mux_module_inst_1_1709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3177]),.i2(intermediate_reg_0[3176]),.o(intermediate_reg_1[1588]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3175]),.i2(intermediate_reg_0[3174]),.o(intermediate_reg_1[1587]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3173]),.i2(intermediate_reg_0[3172]),.o(intermediate_reg_1[1586])); 
mux_module mux_module_inst_1_1712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3171]),.i2(intermediate_reg_0[3170]),.o(intermediate_reg_1[1585]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3169]),.i2(intermediate_reg_0[3168]),.o(intermediate_reg_1[1584]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3167]),.i2(intermediate_reg_0[3166]),.o(intermediate_reg_1[1583])); 
xor_module xor_module_inst_1_1715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3165]),.i2(intermediate_reg_0[3164]),.o(intermediate_reg_1[1582])); 
xor_module xor_module_inst_1_1716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3163]),.i2(intermediate_reg_0[3162]),.o(intermediate_reg_1[1581])); 
xor_module xor_module_inst_1_1717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3161]),.i2(intermediate_reg_0[3160]),.o(intermediate_reg_1[1580])); 
xor_module xor_module_inst_1_1718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3159]),.i2(intermediate_reg_0[3158]),.o(intermediate_reg_1[1579])); 
xor_module xor_module_inst_1_1719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3157]),.i2(intermediate_reg_0[3156]),.o(intermediate_reg_1[1578])); 
xor_module xor_module_inst_1_1720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3155]),.i2(intermediate_reg_0[3154]),.o(intermediate_reg_1[1577])); 
mux_module mux_module_inst_1_1721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3153]),.i2(intermediate_reg_0[3152]),.o(intermediate_reg_1[1576]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3151]),.i2(intermediate_reg_0[3150]),.o(intermediate_reg_1[1575])); 
xor_module xor_module_inst_1_1723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3149]),.i2(intermediate_reg_0[3148]),.o(intermediate_reg_1[1574])); 
mux_module mux_module_inst_1_1724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3147]),.i2(intermediate_reg_0[3146]),.o(intermediate_reg_1[1573]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3145]),.i2(intermediate_reg_0[3144]),.o(intermediate_reg_1[1572])); 
mux_module mux_module_inst_1_1726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3143]),.i2(intermediate_reg_0[3142]),.o(intermediate_reg_1[1571]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3141]),.i2(intermediate_reg_0[3140]),.o(intermediate_reg_1[1570]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3139]),.i2(intermediate_reg_0[3138]),.o(intermediate_reg_1[1569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3137]),.i2(intermediate_reg_0[3136]),.o(intermediate_reg_1[1568]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3135]),.i2(intermediate_reg_0[3134]),.o(intermediate_reg_1[1567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3133]),.i2(intermediate_reg_0[3132]),.o(intermediate_reg_1[1566]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3131]),.i2(intermediate_reg_0[3130]),.o(intermediate_reg_1[1565])); 
xor_module xor_module_inst_1_1733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3129]),.i2(intermediate_reg_0[3128]),.o(intermediate_reg_1[1564])); 
xor_module xor_module_inst_1_1734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3127]),.i2(intermediate_reg_0[3126]),.o(intermediate_reg_1[1563])); 
mux_module mux_module_inst_1_1735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3125]),.i2(intermediate_reg_0[3124]),.o(intermediate_reg_1[1562]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3123]),.i2(intermediate_reg_0[3122]),.o(intermediate_reg_1[1561]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3121]),.i2(intermediate_reg_0[3120]),.o(intermediate_reg_1[1560])); 
mux_module mux_module_inst_1_1738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3119]),.i2(intermediate_reg_0[3118]),.o(intermediate_reg_1[1559]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3117]),.i2(intermediate_reg_0[3116]),.o(intermediate_reg_1[1558])); 
mux_module mux_module_inst_1_1740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3115]),.i2(intermediate_reg_0[3114]),.o(intermediate_reg_1[1557]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3113]),.i2(intermediate_reg_0[3112]),.o(intermediate_reg_1[1556]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3111]),.i2(intermediate_reg_0[3110]),.o(intermediate_reg_1[1555])); 
xor_module xor_module_inst_1_1743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3109]),.i2(intermediate_reg_0[3108]),.o(intermediate_reg_1[1554])); 
mux_module mux_module_inst_1_1744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3107]),.i2(intermediate_reg_0[3106]),.o(intermediate_reg_1[1553]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3105]),.i2(intermediate_reg_0[3104]),.o(intermediate_reg_1[1552])); 
xor_module xor_module_inst_1_1746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3103]),.i2(intermediate_reg_0[3102]),.o(intermediate_reg_1[1551])); 
mux_module mux_module_inst_1_1747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3101]),.i2(intermediate_reg_0[3100]),.o(intermediate_reg_1[1550]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3099]),.i2(intermediate_reg_0[3098]),.o(intermediate_reg_1[1549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3097]),.i2(intermediate_reg_0[3096]),.o(intermediate_reg_1[1548]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3095]),.i2(intermediate_reg_0[3094]),.o(intermediate_reg_1[1547])); 
xor_module xor_module_inst_1_1751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3093]),.i2(intermediate_reg_0[3092]),.o(intermediate_reg_1[1546])); 
mux_module mux_module_inst_1_1752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3091]),.i2(intermediate_reg_0[3090]),.o(intermediate_reg_1[1545]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3089]),.i2(intermediate_reg_0[3088]),.o(intermediate_reg_1[1544])); 
xor_module xor_module_inst_1_1754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3087]),.i2(intermediate_reg_0[3086]),.o(intermediate_reg_1[1543])); 
mux_module mux_module_inst_1_1755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3085]),.i2(intermediate_reg_0[3084]),.o(intermediate_reg_1[1542]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3083]),.i2(intermediate_reg_0[3082]),.o(intermediate_reg_1[1541])); 
mux_module mux_module_inst_1_1757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3081]),.i2(intermediate_reg_0[3080]),.o(intermediate_reg_1[1540]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3079]),.i2(intermediate_reg_0[3078]),.o(intermediate_reg_1[1539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3077]),.i2(intermediate_reg_0[3076]),.o(intermediate_reg_1[1538]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3075]),.i2(intermediate_reg_0[3074]),.o(intermediate_reg_1[1537]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3073]),.i2(intermediate_reg_0[3072]),.o(intermediate_reg_1[1536])); 
xor_module xor_module_inst_1_1762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3071]),.i2(intermediate_reg_0[3070]),.o(intermediate_reg_1[1535])); 
mux_module mux_module_inst_1_1763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3069]),.i2(intermediate_reg_0[3068]),.o(intermediate_reg_1[1534]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3067]),.i2(intermediate_reg_0[3066]),.o(intermediate_reg_1[1533])); 
mux_module mux_module_inst_1_1765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3065]),.i2(intermediate_reg_0[3064]),.o(intermediate_reg_1[1532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3063]),.i2(intermediate_reg_0[3062]),.o(intermediate_reg_1[1531]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3061]),.i2(intermediate_reg_0[3060]),.o(intermediate_reg_1[1530])); 
xor_module xor_module_inst_1_1768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3059]),.i2(intermediate_reg_0[3058]),.o(intermediate_reg_1[1529])); 
mux_module mux_module_inst_1_1769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3057]),.i2(intermediate_reg_0[3056]),.o(intermediate_reg_1[1528]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3055]),.i2(intermediate_reg_0[3054]),.o(intermediate_reg_1[1527]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3053]),.i2(intermediate_reg_0[3052]),.o(intermediate_reg_1[1526])); 
xor_module xor_module_inst_1_1772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3051]),.i2(intermediate_reg_0[3050]),.o(intermediate_reg_1[1525])); 
mux_module mux_module_inst_1_1773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3049]),.i2(intermediate_reg_0[3048]),.o(intermediate_reg_1[1524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3047]),.i2(intermediate_reg_0[3046]),.o(intermediate_reg_1[1523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3045]),.i2(intermediate_reg_0[3044]),.o(intermediate_reg_1[1522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3043]),.i2(intermediate_reg_0[3042]),.o(intermediate_reg_1[1521]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3041]),.i2(intermediate_reg_0[3040]),.o(intermediate_reg_1[1520])); 
xor_module xor_module_inst_1_1778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3039]),.i2(intermediate_reg_0[3038]),.o(intermediate_reg_1[1519])); 
xor_module xor_module_inst_1_1779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3037]),.i2(intermediate_reg_0[3036]),.o(intermediate_reg_1[1518])); 
xor_module xor_module_inst_1_1780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3035]),.i2(intermediate_reg_0[3034]),.o(intermediate_reg_1[1517])); 
xor_module xor_module_inst_1_1781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3033]),.i2(intermediate_reg_0[3032]),.o(intermediate_reg_1[1516])); 
xor_module xor_module_inst_1_1782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3031]),.i2(intermediate_reg_0[3030]),.o(intermediate_reg_1[1515])); 
xor_module xor_module_inst_1_1783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3029]),.i2(intermediate_reg_0[3028]),.o(intermediate_reg_1[1514])); 
mux_module mux_module_inst_1_1784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3027]),.i2(intermediate_reg_0[3026]),.o(intermediate_reg_1[1513]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3025]),.i2(intermediate_reg_0[3024]),.o(intermediate_reg_1[1512])); 
xor_module xor_module_inst_1_1786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3023]),.i2(intermediate_reg_0[3022]),.o(intermediate_reg_1[1511])); 
mux_module mux_module_inst_1_1787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3021]),.i2(intermediate_reg_0[3020]),.o(intermediate_reg_1[1510]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3019]),.i2(intermediate_reg_0[3018]),.o(intermediate_reg_1[1509])); 
xor_module xor_module_inst_1_1789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3017]),.i2(intermediate_reg_0[3016]),.o(intermediate_reg_1[1508])); 
xor_module xor_module_inst_1_1790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3015]),.i2(intermediate_reg_0[3014]),.o(intermediate_reg_1[1507])); 
xor_module xor_module_inst_1_1791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3013]),.i2(intermediate_reg_0[3012]),.o(intermediate_reg_1[1506])); 
xor_module xor_module_inst_1_1792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3011]),.i2(intermediate_reg_0[3010]),.o(intermediate_reg_1[1505])); 
xor_module xor_module_inst_1_1793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3009]),.i2(intermediate_reg_0[3008]),.o(intermediate_reg_1[1504])); 
xor_module xor_module_inst_1_1794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3007]),.i2(intermediate_reg_0[3006]),.o(intermediate_reg_1[1503])); 
xor_module xor_module_inst_1_1795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3005]),.i2(intermediate_reg_0[3004]),.o(intermediate_reg_1[1502])); 
xor_module xor_module_inst_1_1796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3003]),.i2(intermediate_reg_0[3002]),.o(intermediate_reg_1[1501])); 
xor_module xor_module_inst_1_1797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3001]),.i2(intermediate_reg_0[3000]),.o(intermediate_reg_1[1500])); 
mux_module mux_module_inst_1_1798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2999]),.i2(intermediate_reg_0[2998]),.o(intermediate_reg_1[1499]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2997]),.i2(intermediate_reg_0[2996]),.o(intermediate_reg_1[1498]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2995]),.i2(intermediate_reg_0[2994]),.o(intermediate_reg_1[1497])); 
mux_module mux_module_inst_1_1801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2993]),.i2(intermediate_reg_0[2992]),.o(intermediate_reg_1[1496]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2991]),.i2(intermediate_reg_0[2990]),.o(intermediate_reg_1[1495]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2989]),.i2(intermediate_reg_0[2988]),.o(intermediate_reg_1[1494])); 
mux_module mux_module_inst_1_1804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2987]),.i2(intermediate_reg_0[2986]),.o(intermediate_reg_1[1493]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2985]),.i2(intermediate_reg_0[2984]),.o(intermediate_reg_1[1492])); 
mux_module mux_module_inst_1_1806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2983]),.i2(intermediate_reg_0[2982]),.o(intermediate_reg_1[1491]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2981]),.i2(intermediate_reg_0[2980]),.o(intermediate_reg_1[1490])); 
xor_module xor_module_inst_1_1808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2979]),.i2(intermediate_reg_0[2978]),.o(intermediate_reg_1[1489])); 
xor_module xor_module_inst_1_1809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2977]),.i2(intermediate_reg_0[2976]),.o(intermediate_reg_1[1488])); 
mux_module mux_module_inst_1_1810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2975]),.i2(intermediate_reg_0[2974]),.o(intermediate_reg_1[1487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2973]),.i2(intermediate_reg_0[2972]),.o(intermediate_reg_1[1486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2971]),.i2(intermediate_reg_0[2970]),.o(intermediate_reg_1[1485]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2969]),.i2(intermediate_reg_0[2968]),.o(intermediate_reg_1[1484])); 
xor_module xor_module_inst_1_1814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2967]),.i2(intermediate_reg_0[2966]),.o(intermediate_reg_1[1483])); 
xor_module xor_module_inst_1_1815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2965]),.i2(intermediate_reg_0[2964]),.o(intermediate_reg_1[1482])); 
xor_module xor_module_inst_1_1816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2963]),.i2(intermediate_reg_0[2962]),.o(intermediate_reg_1[1481])); 
xor_module xor_module_inst_1_1817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2961]),.i2(intermediate_reg_0[2960]),.o(intermediate_reg_1[1480])); 
xor_module xor_module_inst_1_1818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2959]),.i2(intermediate_reg_0[2958]),.o(intermediate_reg_1[1479])); 
xor_module xor_module_inst_1_1819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2957]),.i2(intermediate_reg_0[2956]),.o(intermediate_reg_1[1478])); 
xor_module xor_module_inst_1_1820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2955]),.i2(intermediate_reg_0[2954]),.o(intermediate_reg_1[1477])); 
xor_module xor_module_inst_1_1821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2953]),.i2(intermediate_reg_0[2952]),.o(intermediate_reg_1[1476])); 
xor_module xor_module_inst_1_1822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2951]),.i2(intermediate_reg_0[2950]),.o(intermediate_reg_1[1475])); 
mux_module mux_module_inst_1_1823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2949]),.i2(intermediate_reg_0[2948]),.o(intermediate_reg_1[1474]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2947]),.i2(intermediate_reg_0[2946]),.o(intermediate_reg_1[1473])); 
mux_module mux_module_inst_1_1825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2945]),.i2(intermediate_reg_0[2944]),.o(intermediate_reg_1[1472]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2943]),.i2(intermediate_reg_0[2942]),.o(intermediate_reg_1[1471])); 
mux_module mux_module_inst_1_1827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2941]),.i2(intermediate_reg_0[2940]),.o(intermediate_reg_1[1470]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2939]),.i2(intermediate_reg_0[2938]),.o(intermediate_reg_1[1469])); 
mux_module mux_module_inst_1_1829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2937]),.i2(intermediate_reg_0[2936]),.o(intermediate_reg_1[1468]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2935]),.i2(intermediate_reg_0[2934]),.o(intermediate_reg_1[1467])); 
mux_module mux_module_inst_1_1831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2933]),.i2(intermediate_reg_0[2932]),.o(intermediate_reg_1[1466]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2931]),.i2(intermediate_reg_0[2930]),.o(intermediate_reg_1[1465])); 
xor_module xor_module_inst_1_1833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2929]),.i2(intermediate_reg_0[2928]),.o(intermediate_reg_1[1464])); 
xor_module xor_module_inst_1_1834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2927]),.i2(intermediate_reg_0[2926]),.o(intermediate_reg_1[1463])); 
mux_module mux_module_inst_1_1835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2925]),.i2(intermediate_reg_0[2924]),.o(intermediate_reg_1[1462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2923]),.i2(intermediate_reg_0[2922]),.o(intermediate_reg_1[1461]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2921]),.i2(intermediate_reg_0[2920]),.o(intermediate_reg_1[1460])); 
mux_module mux_module_inst_1_1838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2919]),.i2(intermediate_reg_0[2918]),.o(intermediate_reg_1[1459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2917]),.i2(intermediate_reg_0[2916]),.o(intermediate_reg_1[1458]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2915]),.i2(intermediate_reg_0[2914]),.o(intermediate_reg_1[1457])); 
xor_module xor_module_inst_1_1841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2913]),.i2(intermediate_reg_0[2912]),.o(intermediate_reg_1[1456])); 
mux_module mux_module_inst_1_1842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2911]),.i2(intermediate_reg_0[2910]),.o(intermediate_reg_1[1455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2909]),.i2(intermediate_reg_0[2908]),.o(intermediate_reg_1[1454]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2907]),.i2(intermediate_reg_0[2906]),.o(intermediate_reg_1[1453])); 
xor_module xor_module_inst_1_1845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2905]),.i2(intermediate_reg_0[2904]),.o(intermediate_reg_1[1452])); 
xor_module xor_module_inst_1_1846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2903]),.i2(intermediate_reg_0[2902]),.o(intermediate_reg_1[1451])); 
mux_module mux_module_inst_1_1847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2901]),.i2(intermediate_reg_0[2900]),.o(intermediate_reg_1[1450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2899]),.i2(intermediate_reg_0[2898]),.o(intermediate_reg_1[1449]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2897]),.i2(intermediate_reg_0[2896]),.o(intermediate_reg_1[1448])); 
xor_module xor_module_inst_1_1850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2895]),.i2(intermediate_reg_0[2894]),.o(intermediate_reg_1[1447])); 
mux_module mux_module_inst_1_1851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2893]),.i2(intermediate_reg_0[2892]),.o(intermediate_reg_1[1446]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2891]),.i2(intermediate_reg_0[2890]),.o(intermediate_reg_1[1445])); 
xor_module xor_module_inst_1_1853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2889]),.i2(intermediate_reg_0[2888]),.o(intermediate_reg_1[1444])); 
mux_module mux_module_inst_1_1854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2887]),.i2(intermediate_reg_0[2886]),.o(intermediate_reg_1[1443]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2885]),.i2(intermediate_reg_0[2884]),.o(intermediate_reg_1[1442]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2883]),.i2(intermediate_reg_0[2882]),.o(intermediate_reg_1[1441])); 
mux_module mux_module_inst_1_1857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2881]),.i2(intermediate_reg_0[2880]),.o(intermediate_reg_1[1440]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2879]),.i2(intermediate_reg_0[2878]),.o(intermediate_reg_1[1439])); 
mux_module mux_module_inst_1_1859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2877]),.i2(intermediate_reg_0[2876]),.o(intermediate_reg_1[1438]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2875]),.i2(intermediate_reg_0[2874]),.o(intermediate_reg_1[1437])); 
mux_module mux_module_inst_1_1861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2873]),.i2(intermediate_reg_0[2872]),.o(intermediate_reg_1[1436]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2871]),.i2(intermediate_reg_0[2870]),.o(intermediate_reg_1[1435])); 
xor_module xor_module_inst_1_1863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2869]),.i2(intermediate_reg_0[2868]),.o(intermediate_reg_1[1434])); 
xor_module xor_module_inst_1_1864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2867]),.i2(intermediate_reg_0[2866]),.o(intermediate_reg_1[1433])); 
xor_module xor_module_inst_1_1865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2865]),.i2(intermediate_reg_0[2864]),.o(intermediate_reg_1[1432])); 
mux_module mux_module_inst_1_1866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2863]),.i2(intermediate_reg_0[2862]),.o(intermediate_reg_1[1431]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2861]),.i2(intermediate_reg_0[2860]),.o(intermediate_reg_1[1430])); 
xor_module xor_module_inst_1_1868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2859]),.i2(intermediate_reg_0[2858]),.o(intermediate_reg_1[1429])); 
xor_module xor_module_inst_1_1869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2857]),.i2(intermediate_reg_0[2856]),.o(intermediate_reg_1[1428])); 
xor_module xor_module_inst_1_1870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2855]),.i2(intermediate_reg_0[2854]),.o(intermediate_reg_1[1427])); 
xor_module xor_module_inst_1_1871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2853]),.i2(intermediate_reg_0[2852]),.o(intermediate_reg_1[1426])); 
mux_module mux_module_inst_1_1872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2851]),.i2(intermediate_reg_0[2850]),.o(intermediate_reg_1[1425]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2849]),.i2(intermediate_reg_0[2848]),.o(intermediate_reg_1[1424]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2847]),.i2(intermediate_reg_0[2846]),.o(intermediate_reg_1[1423]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2845]),.i2(intermediate_reg_0[2844]),.o(intermediate_reg_1[1422])); 
mux_module mux_module_inst_1_1876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2843]),.i2(intermediate_reg_0[2842]),.o(intermediate_reg_1[1421]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2841]),.i2(intermediate_reg_0[2840]),.o(intermediate_reg_1[1420])); 
xor_module xor_module_inst_1_1878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2839]),.i2(intermediate_reg_0[2838]),.o(intermediate_reg_1[1419])); 
xor_module xor_module_inst_1_1879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2837]),.i2(intermediate_reg_0[2836]),.o(intermediate_reg_1[1418])); 
xor_module xor_module_inst_1_1880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2835]),.i2(intermediate_reg_0[2834]),.o(intermediate_reg_1[1417])); 
xor_module xor_module_inst_1_1881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2833]),.i2(intermediate_reg_0[2832]),.o(intermediate_reg_1[1416])); 
xor_module xor_module_inst_1_1882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2831]),.i2(intermediate_reg_0[2830]),.o(intermediate_reg_1[1415])); 
mux_module mux_module_inst_1_1883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2829]),.i2(intermediate_reg_0[2828]),.o(intermediate_reg_1[1414]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2827]),.i2(intermediate_reg_0[2826]),.o(intermediate_reg_1[1413])); 
xor_module xor_module_inst_1_1885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2825]),.i2(intermediate_reg_0[2824]),.o(intermediate_reg_1[1412])); 
xor_module xor_module_inst_1_1886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2823]),.i2(intermediate_reg_0[2822]),.o(intermediate_reg_1[1411])); 
xor_module xor_module_inst_1_1887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2821]),.i2(intermediate_reg_0[2820]),.o(intermediate_reg_1[1410])); 
mux_module mux_module_inst_1_1888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2819]),.i2(intermediate_reg_0[2818]),.o(intermediate_reg_1[1409]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2817]),.i2(intermediate_reg_0[2816]),.o(intermediate_reg_1[1408])); 
xor_module xor_module_inst_1_1890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2815]),.i2(intermediate_reg_0[2814]),.o(intermediate_reg_1[1407])); 
mux_module mux_module_inst_1_1891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2813]),.i2(intermediate_reg_0[2812]),.o(intermediate_reg_1[1406]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2811]),.i2(intermediate_reg_0[2810]),.o(intermediate_reg_1[1405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2809]),.i2(intermediate_reg_0[2808]),.o(intermediate_reg_1[1404]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2807]),.i2(intermediate_reg_0[2806]),.o(intermediate_reg_1[1403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2805]),.i2(intermediate_reg_0[2804]),.o(intermediate_reg_1[1402]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2803]),.i2(intermediate_reg_0[2802]),.o(intermediate_reg_1[1401])); 
xor_module xor_module_inst_1_1897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2801]),.i2(intermediate_reg_0[2800]),.o(intermediate_reg_1[1400])); 
xor_module xor_module_inst_1_1898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2799]),.i2(intermediate_reg_0[2798]),.o(intermediate_reg_1[1399])); 
xor_module xor_module_inst_1_1899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2797]),.i2(intermediate_reg_0[2796]),.o(intermediate_reg_1[1398])); 
mux_module mux_module_inst_1_1900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2795]),.i2(intermediate_reg_0[2794]),.o(intermediate_reg_1[1397]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2793]),.i2(intermediate_reg_0[2792]),.o(intermediate_reg_1[1396])); 
xor_module xor_module_inst_1_1902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2791]),.i2(intermediate_reg_0[2790]),.o(intermediate_reg_1[1395])); 
xor_module xor_module_inst_1_1903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2789]),.i2(intermediate_reg_0[2788]),.o(intermediate_reg_1[1394])); 
xor_module xor_module_inst_1_1904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2787]),.i2(intermediate_reg_0[2786]),.o(intermediate_reg_1[1393])); 
xor_module xor_module_inst_1_1905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2785]),.i2(intermediate_reg_0[2784]),.o(intermediate_reg_1[1392])); 
mux_module mux_module_inst_1_1906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2783]),.i2(intermediate_reg_0[2782]),.o(intermediate_reg_1[1391]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2781]),.i2(intermediate_reg_0[2780]),.o(intermediate_reg_1[1390])); 
mux_module mux_module_inst_1_1908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2779]),.i2(intermediate_reg_0[2778]),.o(intermediate_reg_1[1389]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2777]),.i2(intermediate_reg_0[2776]),.o(intermediate_reg_1[1388]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2775]),.i2(intermediate_reg_0[2774]),.o(intermediate_reg_1[1387])); 
mux_module mux_module_inst_1_1911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2773]),.i2(intermediate_reg_0[2772]),.o(intermediate_reg_1[1386]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2771]),.i2(intermediate_reg_0[2770]),.o(intermediate_reg_1[1385]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2769]),.i2(intermediate_reg_0[2768]),.o(intermediate_reg_1[1384]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2767]),.i2(intermediate_reg_0[2766]),.o(intermediate_reg_1[1383])); 
mux_module mux_module_inst_1_1915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2765]),.i2(intermediate_reg_0[2764]),.o(intermediate_reg_1[1382]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2763]),.i2(intermediate_reg_0[2762]),.o(intermediate_reg_1[1381])); 
mux_module mux_module_inst_1_1917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2761]),.i2(intermediate_reg_0[2760]),.o(intermediate_reg_1[1380]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2759]),.i2(intermediate_reg_0[2758]),.o(intermediate_reg_1[1379]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2757]),.i2(intermediate_reg_0[2756]),.o(intermediate_reg_1[1378])); 
mux_module mux_module_inst_1_1920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2755]),.i2(intermediate_reg_0[2754]),.o(intermediate_reg_1[1377]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2753]),.i2(intermediate_reg_0[2752]),.o(intermediate_reg_1[1376]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2751]),.i2(intermediate_reg_0[2750]),.o(intermediate_reg_1[1375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2749]),.i2(intermediate_reg_0[2748]),.o(intermediate_reg_1[1374]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2747]),.i2(intermediate_reg_0[2746]),.o(intermediate_reg_1[1373]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2745]),.i2(intermediate_reg_0[2744]),.o(intermediate_reg_1[1372])); 
xor_module xor_module_inst_1_1926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2743]),.i2(intermediate_reg_0[2742]),.o(intermediate_reg_1[1371])); 
xor_module xor_module_inst_1_1927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2741]),.i2(intermediate_reg_0[2740]),.o(intermediate_reg_1[1370])); 
mux_module mux_module_inst_1_1928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2739]),.i2(intermediate_reg_0[2738]),.o(intermediate_reg_1[1369]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2737]),.i2(intermediate_reg_0[2736]),.o(intermediate_reg_1[1368])); 
xor_module xor_module_inst_1_1930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2735]),.i2(intermediate_reg_0[2734]),.o(intermediate_reg_1[1367])); 
xor_module xor_module_inst_1_1931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2733]),.i2(intermediate_reg_0[2732]),.o(intermediate_reg_1[1366])); 
mux_module mux_module_inst_1_1932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2731]),.i2(intermediate_reg_0[2730]),.o(intermediate_reg_1[1365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2729]),.i2(intermediate_reg_0[2728]),.o(intermediate_reg_1[1364]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2727]),.i2(intermediate_reg_0[2726]),.o(intermediate_reg_1[1363])); 
mux_module mux_module_inst_1_1935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2725]),.i2(intermediate_reg_0[2724]),.o(intermediate_reg_1[1362]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2723]),.i2(intermediate_reg_0[2722]),.o(intermediate_reg_1[1361])); 
mux_module mux_module_inst_1_1937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2721]),.i2(intermediate_reg_0[2720]),.o(intermediate_reg_1[1360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2719]),.i2(intermediate_reg_0[2718]),.o(intermediate_reg_1[1359]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2717]),.i2(intermediate_reg_0[2716]),.o(intermediate_reg_1[1358])); 
xor_module xor_module_inst_1_1940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2715]),.i2(intermediate_reg_0[2714]),.o(intermediate_reg_1[1357])); 
mux_module mux_module_inst_1_1941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2713]),.i2(intermediate_reg_0[2712]),.o(intermediate_reg_1[1356]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2711]),.i2(intermediate_reg_0[2710]),.o(intermediate_reg_1[1355])); 
mux_module mux_module_inst_1_1943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2709]),.i2(intermediate_reg_0[2708]),.o(intermediate_reg_1[1354]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2707]),.i2(intermediate_reg_0[2706]),.o(intermediate_reg_1[1353])); 
xor_module xor_module_inst_1_1945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2705]),.i2(intermediate_reg_0[2704]),.o(intermediate_reg_1[1352])); 
mux_module mux_module_inst_1_1946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2703]),.i2(intermediate_reg_0[2702]),.o(intermediate_reg_1[1351]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2701]),.i2(intermediate_reg_0[2700]),.o(intermediate_reg_1[1350])); 
mux_module mux_module_inst_1_1948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2699]),.i2(intermediate_reg_0[2698]),.o(intermediate_reg_1[1349]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2697]),.i2(intermediate_reg_0[2696]),.o(intermediate_reg_1[1348]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2695]),.i2(intermediate_reg_0[2694]),.o(intermediate_reg_1[1347]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2693]),.i2(intermediate_reg_0[2692]),.o(intermediate_reg_1[1346]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2691]),.i2(intermediate_reg_0[2690]),.o(intermediate_reg_1[1345]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2689]),.i2(intermediate_reg_0[2688]),.o(intermediate_reg_1[1344])); 
xor_module xor_module_inst_1_1954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2687]),.i2(intermediate_reg_0[2686]),.o(intermediate_reg_1[1343])); 
mux_module mux_module_inst_1_1955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2685]),.i2(intermediate_reg_0[2684]),.o(intermediate_reg_1[1342]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2683]),.i2(intermediate_reg_0[2682]),.o(intermediate_reg_1[1341]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2681]),.i2(intermediate_reg_0[2680]),.o(intermediate_reg_1[1340]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2679]),.i2(intermediate_reg_0[2678]),.o(intermediate_reg_1[1339])); 
mux_module mux_module_inst_1_1959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2677]),.i2(intermediate_reg_0[2676]),.o(intermediate_reg_1[1338]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2675]),.i2(intermediate_reg_0[2674]),.o(intermediate_reg_1[1337]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2673]),.i2(intermediate_reg_0[2672]),.o(intermediate_reg_1[1336])); 
mux_module mux_module_inst_1_1962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2671]),.i2(intermediate_reg_0[2670]),.o(intermediate_reg_1[1335]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2669]),.i2(intermediate_reg_0[2668]),.o(intermediate_reg_1[1334]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2667]),.i2(intermediate_reg_0[2666]),.o(intermediate_reg_1[1333]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2665]),.i2(intermediate_reg_0[2664]),.o(intermediate_reg_1[1332]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2663]),.i2(intermediate_reg_0[2662]),.o(intermediate_reg_1[1331]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2661]),.i2(intermediate_reg_0[2660]),.o(intermediate_reg_1[1330])); 
mux_module mux_module_inst_1_1968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2659]),.i2(intermediate_reg_0[2658]),.o(intermediate_reg_1[1329]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2657]),.i2(intermediate_reg_0[2656]),.o(intermediate_reg_1[1328])); 
xor_module xor_module_inst_1_1970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2655]),.i2(intermediate_reg_0[2654]),.o(intermediate_reg_1[1327])); 
mux_module mux_module_inst_1_1971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2653]),.i2(intermediate_reg_0[2652]),.o(intermediate_reg_1[1326]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2651]),.i2(intermediate_reg_0[2650]),.o(intermediate_reg_1[1325])); 
xor_module xor_module_inst_1_1973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2649]),.i2(intermediate_reg_0[2648]),.o(intermediate_reg_1[1324])); 
mux_module mux_module_inst_1_1974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2647]),.i2(intermediate_reg_0[2646]),.o(intermediate_reg_1[1323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2645]),.i2(intermediate_reg_0[2644]),.o(intermediate_reg_1[1322]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2643]),.i2(intermediate_reg_0[2642]),.o(intermediate_reg_1[1321]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2641]),.i2(intermediate_reg_0[2640]),.o(intermediate_reg_1[1320])); 
xor_module xor_module_inst_1_1978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2639]),.i2(intermediate_reg_0[2638]),.o(intermediate_reg_1[1319])); 
mux_module mux_module_inst_1_1979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2637]),.i2(intermediate_reg_0[2636]),.o(intermediate_reg_1[1318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2635]),.i2(intermediate_reg_0[2634]),.o(intermediate_reg_1[1317]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2633]),.i2(intermediate_reg_0[2632]),.o(intermediate_reg_1[1316])); 
mux_module mux_module_inst_1_1982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2631]),.i2(intermediate_reg_0[2630]),.o(intermediate_reg_1[1315]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2629]),.i2(intermediate_reg_0[2628]),.o(intermediate_reg_1[1314])); 
xor_module xor_module_inst_1_1984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2627]),.i2(intermediate_reg_0[2626]),.o(intermediate_reg_1[1313])); 
xor_module xor_module_inst_1_1985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2625]),.i2(intermediate_reg_0[2624]),.o(intermediate_reg_1[1312])); 
mux_module mux_module_inst_1_1986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309])); 
xor_module xor_module_inst_1_1989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308])); 
xor_module xor_module_inst_1_1990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307])); 
mux_module mux_module_inst_1_1991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303])); 
mux_module mux_module_inst_1_1995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301])); 
xor_module xor_module_inst_1_1997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300])); 
mux_module mux_module_inst_1_1998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297])); 
xor_module xor_module_inst_1_2001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296])); 
mux_module mux_module_inst_1_2002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294])); 
mux_module mux_module_inst_1_2004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290])); 
mux_module mux_module_inst_1_2008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288])); 
mux_module mux_module_inst_1_2010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285])); 
xor_module xor_module_inst_1_2013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284])); 
mux_module mux_module_inst_1_2014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282])); 
mux_module mux_module_inst_1_2016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280])); 
mux_module mux_module_inst_1_2018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276])); 
mux_module mux_module_inst_1_2022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270])); 
mux_module mux_module_inst_1_2028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268])); 
xor_module xor_module_inst_1_2030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267])); 
xor_module xor_module_inst_1_2031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266])); 
xor_module xor_module_inst_1_2032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265])); 
xor_module xor_module_inst_1_2033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264])); 
xor_module xor_module_inst_1_2034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263])); 
xor_module xor_module_inst_1_2035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262])); 
mux_module mux_module_inst_1_2036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257])); 
mux_module mux_module_inst_1_2041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255])); 
mux_module mux_module_inst_1_2043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253])); 
mux_module mux_module_inst_1_2045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249])); 
mux_module mux_module_inst_1_2049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247])); 
xor_module xor_module_inst_1_2051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246])); 
mux_module mux_module_inst_1_2052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244])); 
xor_module xor_module_inst_1_2054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243])); 
xor_module xor_module_inst_1_2055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242])); 
mux_module mux_module_inst_1_2056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240])); 
xor_module xor_module_inst_1_2058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239])); 
xor_module xor_module_inst_1_2059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238])); 
mux_module mux_module_inst_1_2060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234])); 
xor_module xor_module_inst_1_2064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233])); 
xor_module xor_module_inst_1_2065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232])); 
xor_module xor_module_inst_1_2066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231])); 
mux_module mux_module_inst_1_2067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229])); 
mux_module mux_module_inst_1_2069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
mux_module mux_module_inst_1_2072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224])); 
xor_module xor_module_inst_1_2074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223])); 
xor_module xor_module_inst_1_2075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222])); 
xor_module xor_module_inst_1_2076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221])); 
mux_module mux_module_inst_1_2077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218])); 
mux_module mux_module_inst_1_2080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216])); 
mux_module mux_module_inst_1_2082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213])); 
mux_module mux_module_inst_1_2085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210])); 
xor_module xor_module_inst_1_2088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209])); 
mux_module mux_module_inst_1_2089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203])); 
mux_module mux_module_inst_1_2095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201])); 
mux_module mux_module_inst_1_2097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199])); 
mux_module mux_module_inst_1_2099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194])); 
xor_module xor_module_inst_1_2104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193])); 
mux_module mux_module_inst_1_2105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189])); 
mux_module mux_module_inst_1_2109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186])); 
mux_module mux_module_inst_1_2112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184])); 
mux_module mux_module_inst_1_2114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181])); 
xor_module xor_module_inst_1_2117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180])); 
xor_module xor_module_inst_1_2118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179])); 
mux_module mux_module_inst_1_2119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177])); 
mux_module mux_module_inst_1_2121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173])); 
mux_module mux_module_inst_1_2125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167])); 
xor_module xor_module_inst_1_2131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166])); 
mux_module mux_module_inst_1_2132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164])); 
xor_module xor_module_inst_1_2134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163])); 
xor_module xor_module_inst_1_2135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162])); 
xor_module xor_module_inst_1_2136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161])); 
xor_module xor_module_inst_1_2137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160])); 
mux_module mux_module_inst_1_2138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158])); 
xor_module xor_module_inst_1_2140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
xor_module xor_module_inst_1_2141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156])); 
xor_module xor_module_inst_1_2142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155])); 
mux_module mux_module_inst_1_2143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152])); 
mux_module mux_module_inst_1_2146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150])); 
xor_module xor_module_inst_1_2148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149])); 
xor_module xor_module_inst_1_2149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148])); 
xor_module xor_module_inst_1_2150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147])); 
xor_module xor_module_inst_1_2151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146])); 
mux_module mux_module_inst_1_2152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143])); 
xor_module xor_module_inst_1_2155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142])); 
xor_module xor_module_inst_1_2156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141])); 
xor_module xor_module_inst_1_2157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140])); 
mux_module mux_module_inst_1_2158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137])); 
mux_module mux_module_inst_1_2161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135])); 
xor_module xor_module_inst_1_2163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134])); 
mux_module mux_module_inst_1_2164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131])); 
mux_module mux_module_inst_1_2167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127])); 
xor_module xor_module_inst_1_2171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126])); 
xor_module xor_module_inst_1_2172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125])); 
xor_module xor_module_inst_1_2173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124])); 
mux_module mux_module_inst_1_2174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122])); 
mux_module mux_module_inst_1_2176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120])); 
xor_module xor_module_inst_1_2178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119])); 
mux_module mux_module_inst_1_2179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117])); 
mux_module mux_module_inst_1_2181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115])); 
xor_module xor_module_inst_1_2183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114])); 
xor_module xor_module_inst_1_2184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113])); 
xor_module xor_module_inst_1_2185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112])); 
mux_module mux_module_inst_1_2186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110])); 
mux_module mux_module_inst_1_2188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
mux_module mux_module_inst_1_2193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103])); 
xor_module xor_module_inst_1_2195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102])); 
xor_module xor_module_inst_1_2196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
xor_module xor_module_inst_1_2197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100])); 
mux_module mux_module_inst_1_2198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098])); 
mux_module mux_module_inst_1_2200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
xor_module xor_module_inst_1_2205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
xor_module xor_module_inst_1_2206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
mux_module mux_module_inst_1_2207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
xor_module xor_module_inst_1_2209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088])); 
mux_module mux_module_inst_1_2210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
xor_module xor_module_inst_1_2215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082])); 
mux_module mux_module_inst_1_2216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079])); 
mux_module mux_module_inst_1_2219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077])); 
mux_module mux_module_inst_1_2221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075])); 
mux_module mux_module_inst_1_2223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
xor_module xor_module_inst_1_2225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072])); 
xor_module xor_module_inst_1_2226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071])); 
xor_module xor_module_inst_1_2227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070])); 
mux_module mux_module_inst_1_2228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
xor_module xor_module_inst_1_2231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066])); 
xor_module xor_module_inst_1_2232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065])); 
mux_module mux_module_inst_1_2233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062])); 
xor_module xor_module_inst_1_2236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061])); 
xor_module xor_module_inst_1_2237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060])); 
xor_module xor_module_inst_1_2238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059])); 
mux_module mux_module_inst_1_2239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057])); 
mux_module mux_module_inst_1_2241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053])); 
xor_module xor_module_inst_1_2245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
xor_module xor_module_inst_1_2246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051])); 
xor_module xor_module_inst_1_2247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050])); 
xor_module xor_module_inst_1_2248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049])); 
xor_module xor_module_inst_1_2249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048])); 
xor_module xor_module_inst_1_2250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047])); 
mux_module mux_module_inst_1_2251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045])); 
mux_module mux_module_inst_1_2253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
xor_module xor_module_inst_1_2255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
xor_module xor_module_inst_1_2256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041])); 
mux_module mux_module_inst_1_2257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039])); 
xor_module xor_module_inst_1_2259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038])); 
xor_module xor_module_inst_1_2260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037])); 
mux_module mux_module_inst_1_2261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035])); 
xor_module xor_module_inst_1_2263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034])); 
xor_module xor_module_inst_1_2264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033])); 
mux_module mux_module_inst_1_2265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
mux_module mux_module_inst_1_2267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028])); 
xor_module xor_module_inst_1_2270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027])); 
xor_module xor_module_inst_1_2271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026])); 
xor_module xor_module_inst_1_2272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
xor_module xor_module_inst_1_2273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024])); 
xor_module xor_module_inst_1_2274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
xor_module xor_module_inst_1_2275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022])); 
mux_module mux_module_inst_1_2276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
mux_module mux_module_inst_1_2279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
xor_module xor_module_inst_1_2283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
mux_module mux_module_inst_1_2284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012])); 
mux_module mux_module_inst_1_2286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010])); 
xor_module xor_module_inst_1_2288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009])); 
xor_module xor_module_inst_1_2289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
xor_module xor_module_inst_1_2290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
mux_module mux_module_inst_1_2291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
xor_module xor_module_inst_1_2293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004])); 
xor_module xor_module_inst_1_2294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
xor_module xor_module_inst_1_2295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
mux_module mux_module_inst_1_2296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
xor_module xor_module_inst_1_2301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
mux_module mux_module_inst_1_2302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
mux_module mux_module_inst_1_2304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
xor_module xor_module_inst_1_2308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
xor_module xor_module_inst_1_2309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988])); 
mux_module mux_module_inst_1_2310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985])); 
xor_module xor_module_inst_1_2313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
xor_module xor_module_inst_1_2314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
mux_module mux_module_inst_1_2315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
xor_module xor_module_inst_1_2317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
mux_module mux_module_inst_1_2318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
xor_module xor_module_inst_1_2321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
mux_module mux_module_inst_1_2322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974])); 
xor_module xor_module_inst_1_2324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973])); 
xor_module xor_module_inst_1_2325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
mux_module mux_module_inst_1_2326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
xor_module xor_module_inst_1_2329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
mux_module mux_module_inst_1_2330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966])); 
mux_module mux_module_inst_1_2332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
xor_module xor_module_inst_1_2334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
mux_module mux_module_inst_1_2335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
mux_module mux_module_inst_1_2338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
xor_module xor_module_inst_1_2340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957])); 
xor_module xor_module_inst_1_2341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
mux_module mux_module_inst_1_2342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
xor_module xor_module_inst_1_2345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
mux_module mux_module_inst_1_2346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
xor_module xor_module_inst_1_2351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
mux_module mux_module_inst_1_2352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
mux_module mux_module_inst_1_2354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940])); 
mux_module mux_module_inst_1_2358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
xor_module xor_module_inst_1_2363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
mux_module mux_module_inst_1_2364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932])); 
xor_module xor_module_inst_1_2366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
xor_module xor_module_inst_1_2367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930])); 
xor_module xor_module_inst_1_2368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
mux_module mux_module_inst_1_2369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
xor_module xor_module_inst_1_2371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
xor_module xor_module_inst_1_2372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
mux_module mux_module_inst_1_2373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
xor_module xor_module_inst_1_2379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
xor_module xor_module_inst_1_2380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
xor_module xor_module_inst_1_2381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
mux_module mux_module_inst_1_2382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
xor_module xor_module_inst_1_2384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
mux_module mux_module_inst_1_2385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
mux_module mux_module_inst_1_2387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
xor_module xor_module_inst_1_2389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
mux_module mux_module_inst_1_2390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
xor_module xor_module_inst_1_2393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
xor_module xor_module_inst_1_2394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
mux_module mux_module_inst_1_2395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
mux_module mux_module_inst_1_2398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
xor_module xor_module_inst_1_2401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
mux_module mux_module_inst_1_2402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
xor_module xor_module_inst_1_2404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893])); 
xor_module xor_module_inst_1_2405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
xor_module xor_module_inst_1_2406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
xor_module xor_module_inst_1_2407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
mux_module mux_module_inst_1_2408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
mux_module mux_module_inst_1_2410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
xor_module xor_module_inst_1_2415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
xor_module xor_module_inst_1_2416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
xor_module xor_module_inst_1_2417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
mux_module mux_module_inst_1_2418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
mux_module mux_module_inst_1_2420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
xor_module xor_module_inst_1_2423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
mux_module mux_module_inst_1_2424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
mux_module mux_module_inst_1_2426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
mux_module mux_module_inst_1_2428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
mux_module mux_module_inst_1_2430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
mux_module mux_module_inst_1_2432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
mux_module mux_module_inst_1_2435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860])); 
mux_module mux_module_inst_1_2438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856])); 
mux_module mux_module_inst_1_2442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
xor_module xor_module_inst_1_2445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
xor_module xor_module_inst_1_2446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851])); 
mux_module mux_module_inst_1_2447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
mux_module mux_module_inst_1_2449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
mux_module mux_module_inst_1_2451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
xor_module xor_module_inst_1_2460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
xor_module xor_module_inst_1_2461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
mux_module mux_module_inst_1_2462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
mux_module mux_module_inst_1_2466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830])); 
xor_module xor_module_inst_1_2468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829])); 
mux_module mux_module_inst_1_2469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
xor_module xor_module_inst_1_2471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
mux_module mux_module_inst_1_2472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824])); 
mux_module mux_module_inst_1_2474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
mux_module mux_module_inst_1_2479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
xor_module xor_module_inst_1_2481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
xor_module xor_module_inst_1_2482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
xor_module xor_module_inst_1_2483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
mux_module mux_module_inst_1_2484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
mux_module mux_module_inst_1_2487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
mux_module mux_module_inst_1_2492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
xor_module xor_module_inst_1_2496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
xor_module xor_module_inst_1_2497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
mux_module mux_module_inst_1_2498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
mux_module mux_module_inst_1_2500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
xor_module xor_module_inst_1_2504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
mux_module mux_module_inst_1_2505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
xor_module xor_module_inst_1_2508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
xor_module xor_module_inst_1_2509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
mux_module mux_module_inst_1_2510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
mux_module mux_module_inst_1_2513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
xor_module xor_module_inst_1_2516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
mux_module mux_module_inst_1_2517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
mux_module mux_module_inst_1_2519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
mux_module mux_module_inst_1_2524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
xor_module xor_module_inst_1_2531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
mux_module mux_module_inst_1_2532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
xor_module xor_module_inst_1_2535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
mux_module mux_module_inst_1_2536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
xor_module xor_module_inst_1_2543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
mux_module mux_module_inst_1_2544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
mux_module mux_module_inst_1_2547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
mux_module mux_module_inst_1_2550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
xor_module xor_module_inst_1_2554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
mux_module mux_module_inst_1_2555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
mux_module mux_module_inst_1_2558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738])); 
mux_module mux_module_inst_1_2560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
xor_module xor_module_inst_1_2562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
mux_module mux_module_inst_1_2563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
xor_module xor_module_inst_1_2565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
xor_module xor_module_inst_1_2566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
mux_module mux_module_inst_1_2567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
xor_module xor_module_inst_1_2572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
mux_module mux_module_inst_1_2573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
xor_module xor_module_inst_1_2576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
mux_module mux_module_inst_1_2577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
mux_module mux_module_inst_1_2579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
xor_module xor_module_inst_1_2583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
xor_module xor_module_inst_1_2584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
mux_module mux_module_inst_1_2585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
xor_module xor_module_inst_1_2589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
xor_module xor_module_inst_1_2590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
xor_module xor_module_inst_1_2591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
xor_module xor_module_inst_1_2592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
mux_module mux_module_inst_1_2593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
xor_module xor_module_inst_1_2595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
mux_module mux_module_inst_1_2596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
xor_module xor_module_inst_1_2601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
mux_module mux_module_inst_1_2602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
xor_module xor_module_inst_1_2606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
mux_module mux_module_inst_1_2607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
mux_module mux_module_inst_1_2609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
mux_module mux_module_inst_1_2618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
mux_module mux_module_inst_1_2620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
xor_module xor_module_inst_1_2622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
mux_module mux_module_inst_1_2623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
xor_module xor_module_inst_1_2625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
xor_module xor_module_inst_1_2626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_2627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
xor_module xor_module_inst_1_2628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
xor_module xor_module_inst_1_2629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
mux_module mux_module_inst_1_2630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
mux_module mux_module_inst_1_2636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
xor_module xor_module_inst_1_2638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
xor_module xor_module_inst_1_2639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
xor_module xor_module_inst_1_2640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
xor_module xor_module_inst_1_2641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
mux_module mux_module_inst_1_2642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
xor_module xor_module_inst_1_2645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
xor_module xor_module_inst_1_2646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
xor_module xor_module_inst_1_2647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
xor_module xor_module_inst_1_2648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
xor_module xor_module_inst_1_2649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
xor_module xor_module_inst_1_2650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
mux_module mux_module_inst_1_2651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
mux_module mux_module_inst_1_2653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
mux_module mux_module_inst_1_2655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
mux_module mux_module_inst_1_2657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
mux_module mux_module_inst_1_2660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
xor_module xor_module_inst_1_2662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_2663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
mux_module mux_module_inst_1_2664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
mux_module mux_module_inst_1_2672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
mux_module mux_module_inst_1_2674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
xor_module xor_module_inst_1_2677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
mux_module mux_module_inst_1_2678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
xor_module xor_module_inst_1_2680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
mux_module mux_module_inst_1_2681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
xor_module xor_module_inst_1_2683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
xor_module xor_module_inst_1_2684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
xor_module xor_module_inst_1_2685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
mux_module mux_module_inst_1_2686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
mux_module mux_module_inst_1_2689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
mux_module mux_module_inst_1_2693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
mux_module mux_module_inst_1_2698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
mux_module mux_module_inst_1_2700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
xor_module xor_module_inst_1_2702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
mux_module mux_module_inst_1_2703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
mux_module mux_module_inst_1_2705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
xor_module xor_module_inst_1_2710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
xor_module xor_module_inst_1_2711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
mux_module mux_module_inst_1_2712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
mux_module mux_module_inst_1_2714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
xor_module xor_module_inst_1_2716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
mux_module mux_module_inst_1_2717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
xor_module xor_module_inst_1_2720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
xor_module xor_module_inst_1_2721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
xor_module xor_module_inst_1_2722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
mux_module mux_module_inst_1_2723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
xor_module xor_module_inst_1_2727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
xor_module xor_module_inst_1_2728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
mux_module mux_module_inst_1_2729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
xor_module xor_module_inst_1_2734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
mux_module mux_module_inst_1_2735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
xor_module xor_module_inst_1_2737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
mux_module mux_module_inst_1_2738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
xor_module xor_module_inst_1_2742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
mux_module mux_module_inst_1_2743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
xor_module xor_module_inst_1_2745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
xor_module xor_module_inst_1_2746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
xor_module xor_module_inst_1_2747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
mux_module mux_module_inst_1_2748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
mux_module mux_module_inst_1_2751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
xor_module xor_module_inst_1_2753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
xor_module xor_module_inst_1_2754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
xor_module xor_module_inst_1_2755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
xor_module xor_module_inst_1_2756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
mux_module mux_module_inst_1_2757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
mux_module mux_module_inst_1_2759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
xor_module xor_module_inst_1_2762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
mux_module mux_module_inst_1_2763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
mux_module mux_module_inst_1_2766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
mux_module mux_module_inst_1_2768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
mux_module mux_module_inst_1_2772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
xor_module xor_module_inst_1_2783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
xor_module xor_module_inst_1_2784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
xor_module xor_module_inst_1_2785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
mux_module mux_module_inst_1_2786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
mux_module mux_module_inst_1_2788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
xor_module xor_module_inst_1_2790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
xor_module xor_module_inst_1_2791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
xor_module xor_module_inst_1_2792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
xor_module xor_module_inst_1_2793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
mux_module mux_module_inst_1_2794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
xor_module xor_module_inst_1_2802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
xor_module xor_module_inst_1_2803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
mux_module mux_module_inst_1_2804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
mux_module mux_module_inst_1_2807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
mux_module mux_module_inst_1_2809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
xor_module xor_module_inst_1_2812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
xor_module xor_module_inst_1_2813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
xor_module xor_module_inst_1_2814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
xor_module xor_module_inst_1_2815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_2816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
mux_module mux_module_inst_1_2818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
xor_module xor_module_inst_1_2821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
xor_module xor_module_inst_1_2822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
mux_module mux_module_inst_1_2823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
xor_module xor_module_inst_1_2826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
xor_module xor_module_inst_1_2827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
xor_module xor_module_inst_1_2828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
mux_module mux_module_inst_1_2829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
xor_module xor_module_inst_1_2831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
xor_module xor_module_inst_1_2832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
xor_module xor_module_inst_1_2833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
mux_module mux_module_inst_1_2834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
mux_module mux_module_inst_1_2838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
xor_module xor_module_inst_1_2841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
xor_module xor_module_inst_1_2842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
mux_module mux_module_inst_1_2843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
mux_module mux_module_inst_1_2847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
mux_module mux_module_inst_1_2849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
xor_module xor_module_inst_1_2851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
xor_module xor_module_inst_1_2852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
xor_module xor_module_inst_1_2853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
mux_module mux_module_inst_1_2854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
xor_module xor_module_inst_1_2856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
mux_module mux_module_inst_1_2857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
mux_module mux_module_inst_1_2862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
mux_module mux_module_inst_1_2866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
mux_module mux_module_inst_1_2871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
xor_module xor_module_inst_1_2873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
mux_module mux_module_inst_1_2874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
mux_module mux_module_inst_1_2876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
mux_module mux_module_inst_1_2879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
xor_module xor_module_inst_1_2881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
xor_module xor_module_inst_1_2882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
mux_module mux_module_inst_1_2883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
xor_module xor_module_inst_1_2889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
xor_module xor_module_inst_1_2890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
mux_module mux_module_inst_1_2891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
xor_module xor_module_inst_1_2893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
xor_module xor_module_inst_1_2894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
mux_module mux_module_inst_1_2895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
mux_module mux_module_inst_1_2897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
mux_module mux_module_inst_1_2899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
mux_module mux_module_inst_1_2901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
mux_module mux_module_inst_1_2903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
xor_module xor_module_inst_1_2905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
xor_module xor_module_inst_1_2906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
xor_module xor_module_inst_1_2907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_2908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
mux_module mux_module_inst_1_2909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
mux_module mux_module_inst_1_2911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
xor_module xor_module_inst_1_2914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
mux_module mux_module_inst_1_2915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
xor_module xor_module_inst_1_2918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
mux_module mux_module_inst_1_2919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
xor_module xor_module_inst_1_2921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_2922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
xor_module xor_module_inst_1_2927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
xor_module xor_module_inst_1_2928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
mux_module mux_module_inst_1_2929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
xor_module xor_module_inst_1_2931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
xor_module xor_module_inst_1_2932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
mux_module mux_module_inst_1_2933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
mux_module mux_module_inst_1_2935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
mux_module mux_module_inst_1_2937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
mux_module mux_module_inst_1_2939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
mux_module mux_module_inst_1_2941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
xor_module xor_module_inst_1_2946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
mux_module mux_module_inst_1_2947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
xor_module xor_module_inst_1_2949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
xor_module xor_module_inst_1_2950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
xor_module xor_module_inst_1_2951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
xor_module xor_module_inst_1_2952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
xor_module xor_module_inst_1_2953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
xor_module xor_module_inst_1_2954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
xor_module xor_module_inst_1_2955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
xor_module xor_module_inst_1_2956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
mux_module mux_module_inst_1_2957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
mux_module mux_module_inst_1_2959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
xor_module xor_module_inst_1_2961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
xor_module xor_module_inst_1_2962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
xor_module xor_module_inst_1_2963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
xor_module xor_module_inst_1_2964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
mux_module mux_module_inst_1_2965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
mux_module mux_module_inst_1_2968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
xor_module xor_module_inst_1_2970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
mux_module mux_module_inst_1_2971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
mux_module mux_module_inst_1_2974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
mux_module mux_module_inst_1_2977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
xor_module xor_module_inst_1_2981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
mux_module mux_module_inst_1_2982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
xor_module xor_module_inst_1_2985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
xor_module xor_module_inst_1_2986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
mux_module mux_module_inst_1_2987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
mux_module mux_module_inst_1_2990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
mux_module mux_module_inst_1_2993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
xor_module xor_module_inst_1_2997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
xor_module xor_module_inst_1_2998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
xor_module xor_module_inst_1_2999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
mux_module mux_module_inst_1_3000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
mux_module mux_module_inst_1_3002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
mux_module mux_module_inst_1_3004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
xor_module xor_module_inst_1_3006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
xor_module xor_module_inst_1_3007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
xor_module xor_module_inst_1_3008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_3009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
mux_module mux_module_inst_1_3010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
xor_module xor_module_inst_1_3012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
mux_module mux_module_inst_1_3013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
mux_module mux_module_inst_1_3016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
xor_module xor_module_inst_1_3018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
xor_module xor_module_inst_1_3019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
mux_module mux_module_inst_1_3020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
xor_module xor_module_inst_1_3027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
xor_module xor_module_inst_1_3028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
xor_module xor_module_inst_1_3029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
xor_module xor_module_inst_1_3030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
xor_module xor_module_inst_1_3031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
mux_module mux_module_inst_1_3032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
xor_module xor_module_inst_1_3034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
mux_module mux_module_inst_1_3035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
xor_module xor_module_inst_1_3037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
mux_module mux_module_inst_1_3038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
mux_module mux_module_inst_1_3040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
mux_module mux_module_inst_1_3042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
xor_module xor_module_inst_1_3045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
mux_module mux_module_inst_1_3046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
xor_module xor_module_inst_1_3048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
xor_module xor_module_inst_1_3049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
xor_module xor_module_inst_1_3050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
xor_module xor_module_inst_1_3051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
mux_module mux_module_inst_1_3052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
xor_module xor_module_inst_1_3055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
xor_module xor_module_inst_1_3056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
mux_module mux_module_inst_1_3057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
mux_module mux_module_inst_1_3061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
mux_module mux_module_inst_1_3064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
xor_module xor_module_inst_1_3067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_3068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
xor_module xor_module_inst_1_3069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
xor_module xor_module_inst_1_3070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
mux_module mux_module_inst_1_3071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
mux_module mux_module_inst_1_3076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
xor_module xor_module_inst_1_3079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
mux_module mux_module_inst_1_3080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
xor_module xor_module_inst_1_3083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
xor_module xor_module_inst_1_3084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
xor_module xor_module_inst_1_3085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
mux_module mux_module_inst_1_3086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
xor_module xor_module_inst_1_3090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
xor_module xor_module_inst_1_3091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
xor_module xor_module_inst_1_3092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
mux_module mux_module_inst_1_3093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
mux_module mux_module_inst_1_3101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
mux_module mux_module_inst_1_3103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
mux_module mux_module_inst_1_3106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
xor_module xor_module_inst_1_3108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
xor_module xor_module_inst_1_3109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
xor_module xor_module_inst_1_3110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
mux_module mux_module_inst_1_3111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
mux_module mux_module_inst_1_3113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
xor_module xor_module_inst_1_3115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
xor_module xor_module_inst_1_3116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
mux_module mux_module_inst_1_3117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
mux_module mux_module_inst_1_3120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
xor_module xor_module_inst_1_3122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
xor_module xor_module_inst_1_3123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
xor_module xor_module_inst_1_3124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
mux_module mux_module_inst_1_3125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
xor_module xor_module_inst_1_3128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
mux_module mux_module_inst_1_3129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
mux_module mux_module_inst_1_3131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
mux_module mux_module_inst_1_3133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
xor_module xor_module_inst_1_3136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
xor_module xor_module_inst_1_3137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
mux_module mux_module_inst_1_3138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
mux_module mux_module_inst_1_3140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_3143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
mux_module mux_module_inst_1_3144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
mux_module mux_module_inst_1_3146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
mux_module mux_module_inst_1_3149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
mux_module mux_module_inst_1_3151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
mux_module mux_module_inst_1_3153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
mux_module mux_module_inst_1_3160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
xor_module xor_module_inst_1_3165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
mux_module mux_module_inst_1_3166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
mux_module mux_module_inst_1_3168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
xor_module xor_module_inst_1_3170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
mux_module mux_module_inst_1_3171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
xor_module xor_module_inst_1_3174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
xor_module xor_module_inst_1_3175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
xor_module xor_module_inst_1_3176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
xor_module xor_module_inst_1_3177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
mux_module mux_module_inst_1_3178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
xor_module xor_module_inst_1_3181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
xor_module xor_module_inst_1_3182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
xor_module xor_module_inst_1_3183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
xor_module xor_module_inst_1_3184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
xor_module xor_module_inst_1_3185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
mux_module mux_module_inst_1_3186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
xor_module xor_module_inst_1_3188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
xor_module xor_module_inst_1_3189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
xor_module xor_module_inst_1_3190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
mux_module mux_module_inst_1_3191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
xor_module xor_module_inst_1_3193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
xor_module xor_module_inst_1_3194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
xor_module xor_module_inst_1_3195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
xor_module xor_module_inst_1_3196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
mux_module mux_module_inst_1_3197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
xor_module xor_module_inst_1_3199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
xor_module xor_module_inst_1_3200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
mux_module mux_module_inst_1_3201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
xor_module xor_module_inst_1_3203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
mux_module mux_module_inst_1_3204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
xor_module xor_module_inst_1_3206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
xor_module xor_module_inst_1_3207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
xor_module xor_module_inst_1_3208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
mux_module mux_module_inst_1_3209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
xor_module xor_module_inst_1_3211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
xor_module xor_module_inst_1_3212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
mux_module mux_module_inst_1_3213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
mux_module mux_module_inst_1_3215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
mux_module mux_module_inst_1_3219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
mux_module mux_module_inst_1_3221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
xor_module xor_module_inst_1_3224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
xor_module xor_module_inst_1_3225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
mux_module mux_module_inst_1_3226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
mux_module mux_module_inst_1_3228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
mux_module mux_module_inst_1_3231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
mux_module mux_module_inst_1_3234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
xor_module xor_module_inst_1_3239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
mux_module mux_module_inst_1_3240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
mux_module mux_module_inst_1_3242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
mux_module mux_module_inst_1_3245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
xor_module xor_module_inst_1_3247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
mux_module mux_module_inst_1_3248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
xor_module xor_module_inst_1_3251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
xor_module xor_module_inst_1_3252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
mux_module mux_module_inst_1_3253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
mux_module mux_module_inst_1_3256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
mux_module mux_module_inst_1_3258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
mux_module mux_module_inst_1_3264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
xor_module xor_module_inst_1_3266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
mux_module mux_module_inst_1_3267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
mux_module mux_module_inst_1_3271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
xor_module xor_module_inst_1_3273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
mux_module mux_module_inst_1_3274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
mux_module mux_module_inst_1_3278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
xor_module xor_module_inst_1_3282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
xor_module xor_module_inst_1_3283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
mux_module mux_module_inst_1_3284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
xor_module xor_module_inst_1_3286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
xor_module xor_module_inst_1_3287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
mux_module mux_module_inst_1_3288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
xor_module xor_module_inst_1_3290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
mux_module mux_module_inst_1_3291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
xor_module xor_module_inst_1_3295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
mux_module mux_module_inst_1_3296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
wire [1648:0]intermediate_reg_2; 
 
xor_module xor_module_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3297]),.i2(intermediate_reg_1[3296]),.o(intermediate_reg_2[1648])); 
mux_module mux_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3295]),.i2(intermediate_reg_1[3294]),.o(intermediate_reg_2[1647]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3293]),.i2(intermediate_reg_1[3292]),.o(intermediate_reg_2[1646]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3291]),.i2(intermediate_reg_1[3290]),.o(intermediate_reg_2[1645]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3289]),.i2(intermediate_reg_1[3288]),.o(intermediate_reg_2[1644]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3287]),.i2(intermediate_reg_1[3286]),.o(intermediate_reg_2[1643]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3285]),.i2(intermediate_reg_1[3284]),.o(intermediate_reg_2[1642]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3283]),.i2(intermediate_reg_1[3282]),.o(intermediate_reg_2[1641]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3281]),.i2(intermediate_reg_1[3280]),.o(intermediate_reg_2[1640]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3279]),.i2(intermediate_reg_1[3278]),.o(intermediate_reg_2[1639]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3277]),.i2(intermediate_reg_1[3276]),.o(intermediate_reg_2[1638])); 
mux_module mux_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3275]),.i2(intermediate_reg_1[3274]),.o(intermediate_reg_2[1637]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3273]),.i2(intermediate_reg_1[3272]),.o(intermediate_reg_2[1636]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3271]),.i2(intermediate_reg_1[3270]),.o(intermediate_reg_2[1635]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3269]),.i2(intermediate_reg_1[3268]),.o(intermediate_reg_2[1634])); 
mux_module mux_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3267]),.i2(intermediate_reg_1[3266]),.o(intermediate_reg_2[1633]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3265]),.i2(intermediate_reg_1[3264]),.o(intermediate_reg_2[1632]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3263]),.i2(intermediate_reg_1[3262]),.o(intermediate_reg_2[1631]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3261]),.i2(intermediate_reg_1[3260]),.o(intermediate_reg_2[1630])); 
xor_module xor_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3259]),.i2(intermediate_reg_1[3258]),.o(intermediate_reg_2[1629])); 
xor_module xor_module_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3257]),.i2(intermediate_reg_1[3256]),.o(intermediate_reg_2[1628])); 
mux_module mux_module_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3255]),.i2(intermediate_reg_1[3254]),.o(intermediate_reg_2[1627]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3253]),.i2(intermediate_reg_1[3252]),.o(intermediate_reg_2[1626]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3251]),.i2(intermediate_reg_1[3250]),.o(intermediate_reg_2[1625]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3249]),.i2(intermediate_reg_1[3248]),.o(intermediate_reg_2[1624]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3247]),.i2(intermediate_reg_1[3246]),.o(intermediate_reg_2[1623]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3245]),.i2(intermediate_reg_1[3244]),.o(intermediate_reg_2[1622]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3243]),.i2(intermediate_reg_1[3242]),.o(intermediate_reg_2[1621])); 
xor_module xor_module_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3241]),.i2(intermediate_reg_1[3240]),.o(intermediate_reg_2[1620])); 
xor_module xor_module_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3239]),.i2(intermediate_reg_1[3238]),.o(intermediate_reg_2[1619])); 
xor_module xor_module_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3237]),.i2(intermediate_reg_1[3236]),.o(intermediate_reg_2[1618])); 
xor_module xor_module_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3235]),.i2(intermediate_reg_1[3234]),.o(intermediate_reg_2[1617])); 
xor_module xor_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3233]),.i2(intermediate_reg_1[3232]),.o(intermediate_reg_2[1616])); 
mux_module mux_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3231]),.i2(intermediate_reg_1[3230]),.o(intermediate_reg_2[1615]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3229]),.i2(intermediate_reg_1[3228]),.o(intermediate_reg_2[1614])); 
xor_module xor_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3227]),.i2(intermediate_reg_1[3226]),.o(intermediate_reg_2[1613])); 
xor_module xor_module_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3225]),.i2(intermediate_reg_1[3224]),.o(intermediate_reg_2[1612])); 
xor_module xor_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3223]),.i2(intermediate_reg_1[3222]),.o(intermediate_reg_2[1611])); 
xor_module xor_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3221]),.i2(intermediate_reg_1[3220]),.o(intermediate_reg_2[1610])); 
mux_module mux_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3219]),.i2(intermediate_reg_1[3218]),.o(intermediate_reg_2[1609]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3217]),.i2(intermediate_reg_1[3216]),.o(intermediate_reg_2[1608])); 
mux_module mux_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3215]),.i2(intermediate_reg_1[3214]),.o(intermediate_reg_2[1607]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3213]),.i2(intermediate_reg_1[3212]),.o(intermediate_reg_2[1606]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3211]),.i2(intermediate_reg_1[3210]),.o(intermediate_reg_2[1605])); 
xor_module xor_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3209]),.i2(intermediate_reg_1[3208]),.o(intermediate_reg_2[1604])); 
mux_module mux_module_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3207]),.i2(intermediate_reg_1[3206]),.o(intermediate_reg_2[1603]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3205]),.i2(intermediate_reg_1[3204]),.o(intermediate_reg_2[1602])); 
mux_module mux_module_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3203]),.i2(intermediate_reg_1[3202]),.o(intermediate_reg_2[1601]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3201]),.i2(intermediate_reg_1[3200]),.o(intermediate_reg_2[1600])); 
xor_module xor_module_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3199]),.i2(intermediate_reg_1[3198]),.o(intermediate_reg_2[1599])); 
xor_module xor_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3197]),.i2(intermediate_reg_1[3196]),.o(intermediate_reg_2[1598])); 
mux_module mux_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3195]),.i2(intermediate_reg_1[3194]),.o(intermediate_reg_2[1597]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3193]),.i2(intermediate_reg_1[3192]),.o(intermediate_reg_2[1596])); 
xor_module xor_module_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3191]),.i2(intermediate_reg_1[3190]),.o(intermediate_reg_2[1595])); 
xor_module xor_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3189]),.i2(intermediate_reg_1[3188]),.o(intermediate_reg_2[1594])); 
xor_module xor_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3187]),.i2(intermediate_reg_1[3186]),.o(intermediate_reg_2[1593])); 
xor_module xor_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3185]),.i2(intermediate_reg_1[3184]),.o(intermediate_reg_2[1592])); 
mux_module mux_module_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3183]),.i2(intermediate_reg_1[3182]),.o(intermediate_reg_2[1591]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3181]),.i2(intermediate_reg_1[3180]),.o(intermediate_reg_2[1590])); 
xor_module xor_module_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3179]),.i2(intermediate_reg_1[3178]),.o(intermediate_reg_2[1589])); 
mux_module mux_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3177]),.i2(intermediate_reg_1[3176]),.o(intermediate_reg_2[1588]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3175]),.i2(intermediate_reg_1[3174]),.o(intermediate_reg_2[1587])); 
mux_module mux_module_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3173]),.i2(intermediate_reg_1[3172]),.o(intermediate_reg_2[1586]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3171]),.i2(intermediate_reg_1[3170]),.o(intermediate_reg_2[1585]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3169]),.i2(intermediate_reg_1[3168]),.o(intermediate_reg_2[1584]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3167]),.i2(intermediate_reg_1[3166]),.o(intermediate_reg_2[1583])); 
xor_module xor_module_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3165]),.i2(intermediate_reg_1[3164]),.o(intermediate_reg_2[1582])); 
xor_module xor_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3163]),.i2(intermediate_reg_1[3162]),.o(intermediate_reg_2[1581])); 
xor_module xor_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3161]),.i2(intermediate_reg_1[3160]),.o(intermediate_reg_2[1580])); 
xor_module xor_module_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3159]),.i2(intermediate_reg_1[3158]),.o(intermediate_reg_2[1579])); 
xor_module xor_module_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3157]),.i2(intermediate_reg_1[3156]),.o(intermediate_reg_2[1578])); 
xor_module xor_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3155]),.i2(intermediate_reg_1[3154]),.o(intermediate_reg_2[1577])); 
mux_module mux_module_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3153]),.i2(intermediate_reg_1[3152]),.o(intermediate_reg_2[1576]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3151]),.i2(intermediate_reg_1[3150]),.o(intermediate_reg_2[1575]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3149]),.i2(intermediate_reg_1[3148]),.o(intermediate_reg_2[1574])); 
mux_module mux_module_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3147]),.i2(intermediate_reg_1[3146]),.o(intermediate_reg_2[1573]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3145]),.i2(intermediate_reg_1[3144]),.o(intermediate_reg_2[1572]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3143]),.i2(intermediate_reg_1[3142]),.o(intermediate_reg_2[1571])); 
xor_module xor_module_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3141]),.i2(intermediate_reg_1[3140]),.o(intermediate_reg_2[1570])); 
mux_module mux_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3139]),.i2(intermediate_reg_1[3138]),.o(intermediate_reg_2[1569]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3137]),.i2(intermediate_reg_1[3136]),.o(intermediate_reg_2[1568])); 
mux_module mux_module_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3135]),.i2(intermediate_reg_1[3134]),.o(intermediate_reg_2[1567]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3133]),.i2(intermediate_reg_1[3132]),.o(intermediate_reg_2[1566]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3131]),.i2(intermediate_reg_1[3130]),.o(intermediate_reg_2[1565]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3129]),.i2(intermediate_reg_1[3128]),.o(intermediate_reg_2[1564]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3127]),.i2(intermediate_reg_1[3126]),.o(intermediate_reg_2[1563])); 
mux_module mux_module_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3125]),.i2(intermediate_reg_1[3124]),.o(intermediate_reg_2[1562]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3123]),.i2(intermediate_reg_1[3122]),.o(intermediate_reg_2[1561]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3121]),.i2(intermediate_reg_1[3120]),.o(intermediate_reg_2[1560]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3119]),.i2(intermediate_reg_1[3118]),.o(intermediate_reg_2[1559])); 
mux_module mux_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3117]),.i2(intermediate_reg_1[3116]),.o(intermediate_reg_2[1558]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3115]),.i2(intermediate_reg_1[3114]),.o(intermediate_reg_2[1557]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3113]),.i2(intermediate_reg_1[3112]),.o(intermediate_reg_2[1556]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3111]),.i2(intermediate_reg_1[3110]),.o(intermediate_reg_2[1555]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3109]),.i2(intermediate_reg_1[3108]),.o(intermediate_reg_2[1554])); 
mux_module mux_module_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3107]),.i2(intermediate_reg_1[3106]),.o(intermediate_reg_2[1553]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3105]),.i2(intermediate_reg_1[3104]),.o(intermediate_reg_2[1552])); 
mux_module mux_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3103]),.i2(intermediate_reg_1[3102]),.o(intermediate_reg_2[1551]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3101]),.i2(intermediate_reg_1[3100]),.o(intermediate_reg_2[1550]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3099]),.i2(intermediate_reg_1[3098]),.o(intermediate_reg_2[1549])); 
mux_module mux_module_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3097]),.i2(intermediate_reg_1[3096]),.o(intermediate_reg_2[1548]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3095]),.i2(intermediate_reg_1[3094]),.o(intermediate_reg_2[1547]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3093]),.i2(intermediate_reg_1[3092]),.o(intermediate_reg_2[1546])); 
mux_module mux_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3091]),.i2(intermediate_reg_1[3090]),.o(intermediate_reg_2[1545]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3089]),.i2(intermediate_reg_1[3088]),.o(intermediate_reg_2[1544]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3087]),.i2(intermediate_reg_1[3086]),.o(intermediate_reg_2[1543]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3085]),.i2(intermediate_reg_1[3084]),.o(intermediate_reg_2[1542]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3083]),.i2(intermediate_reg_1[3082]),.o(intermediate_reg_2[1541])); 
xor_module xor_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3081]),.i2(intermediate_reg_1[3080]),.o(intermediate_reg_2[1540])); 
xor_module xor_module_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3079]),.i2(intermediate_reg_1[3078]),.o(intermediate_reg_2[1539])); 
mux_module mux_module_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3077]),.i2(intermediate_reg_1[3076]),.o(intermediate_reg_2[1538]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3075]),.i2(intermediate_reg_1[3074]),.o(intermediate_reg_2[1537])); 
xor_module xor_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3073]),.i2(intermediate_reg_1[3072]),.o(intermediate_reg_2[1536])); 
xor_module xor_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3071]),.i2(intermediate_reg_1[3070]),.o(intermediate_reg_2[1535])); 
mux_module mux_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3069]),.i2(intermediate_reg_1[3068]),.o(intermediate_reg_2[1534]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3067]),.i2(intermediate_reg_1[3066]),.o(intermediate_reg_2[1533])); 
xor_module xor_module_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3065]),.i2(intermediate_reg_1[3064]),.o(intermediate_reg_2[1532])); 
xor_module xor_module_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3063]),.i2(intermediate_reg_1[3062]),.o(intermediate_reg_2[1531])); 
mux_module mux_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3061]),.i2(intermediate_reg_1[3060]),.o(intermediate_reg_2[1530]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3059]),.i2(intermediate_reg_1[3058]),.o(intermediate_reg_2[1529])); 
xor_module xor_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3057]),.i2(intermediate_reg_1[3056]),.o(intermediate_reg_2[1528])); 
mux_module mux_module_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3055]),.i2(intermediate_reg_1[3054]),.o(intermediate_reg_2[1527]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3053]),.i2(intermediate_reg_1[3052]),.o(intermediate_reg_2[1526]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3051]),.i2(intermediate_reg_1[3050]),.o(intermediate_reg_2[1525])); 
xor_module xor_module_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3049]),.i2(intermediate_reg_1[3048]),.o(intermediate_reg_2[1524])); 
xor_module xor_module_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3047]),.i2(intermediate_reg_1[3046]),.o(intermediate_reg_2[1523])); 
xor_module xor_module_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3045]),.i2(intermediate_reg_1[3044]),.o(intermediate_reg_2[1522])); 
xor_module xor_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3043]),.i2(intermediate_reg_1[3042]),.o(intermediate_reg_2[1521])); 
xor_module xor_module_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3041]),.i2(intermediate_reg_1[3040]),.o(intermediate_reg_2[1520])); 
mux_module mux_module_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3039]),.i2(intermediate_reg_1[3038]),.o(intermediate_reg_2[1519]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3037]),.i2(intermediate_reg_1[3036]),.o(intermediate_reg_2[1518]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3035]),.i2(intermediate_reg_1[3034]),.o(intermediate_reg_2[1517])); 
xor_module xor_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3033]),.i2(intermediate_reg_1[3032]),.o(intermediate_reg_2[1516])); 
mux_module mux_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3031]),.i2(intermediate_reg_1[3030]),.o(intermediate_reg_2[1515]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3029]),.i2(intermediate_reg_1[3028]),.o(intermediate_reg_2[1514]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3027]),.i2(intermediate_reg_1[3026]),.o(intermediate_reg_2[1513])); 
xor_module xor_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3025]),.i2(intermediate_reg_1[3024]),.o(intermediate_reg_2[1512])); 
xor_module xor_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3023]),.i2(intermediate_reg_1[3022]),.o(intermediate_reg_2[1511])); 
mux_module mux_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3021]),.i2(intermediate_reg_1[3020]),.o(intermediate_reg_2[1510]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3019]),.i2(intermediate_reg_1[3018]),.o(intermediate_reg_2[1509]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3017]),.i2(intermediate_reg_1[3016]),.o(intermediate_reg_2[1508])); 
mux_module mux_module_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3015]),.i2(intermediate_reg_1[3014]),.o(intermediate_reg_2[1507]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3013]),.i2(intermediate_reg_1[3012]),.o(intermediate_reg_2[1506])); 
mux_module mux_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3011]),.i2(intermediate_reg_1[3010]),.o(intermediate_reg_2[1505]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3009]),.i2(intermediate_reg_1[3008]),.o(intermediate_reg_2[1504])); 
xor_module xor_module_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3007]),.i2(intermediate_reg_1[3006]),.o(intermediate_reg_2[1503])); 
xor_module xor_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3005]),.i2(intermediate_reg_1[3004]),.o(intermediate_reg_2[1502])); 
xor_module xor_module_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3003]),.i2(intermediate_reg_1[3002]),.o(intermediate_reg_2[1501])); 
mux_module mux_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3001]),.i2(intermediate_reg_1[3000]),.o(intermediate_reg_2[1500]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2999]),.i2(intermediate_reg_1[2998]),.o(intermediate_reg_2[1499])); 
xor_module xor_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2997]),.i2(intermediate_reg_1[2996]),.o(intermediate_reg_2[1498])); 
mux_module mux_module_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2995]),.i2(intermediate_reg_1[2994]),.o(intermediate_reg_2[1497]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2993]),.i2(intermediate_reg_1[2992]),.o(intermediate_reg_2[1496]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2991]),.i2(intermediate_reg_1[2990]),.o(intermediate_reg_2[1495]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2989]),.i2(intermediate_reg_1[2988]),.o(intermediate_reg_2[1494])); 
mux_module mux_module_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2987]),.i2(intermediate_reg_1[2986]),.o(intermediate_reg_2[1493]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2985]),.i2(intermediate_reg_1[2984]),.o(intermediate_reg_2[1492]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2983]),.i2(intermediate_reg_1[2982]),.o(intermediate_reg_2[1491])); 
xor_module xor_module_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2981]),.i2(intermediate_reg_1[2980]),.o(intermediate_reg_2[1490])); 
mux_module mux_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2979]),.i2(intermediate_reg_1[2978]),.o(intermediate_reg_2[1489]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2977]),.i2(intermediate_reg_1[2976]),.o(intermediate_reg_2[1488])); 
xor_module xor_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2975]),.i2(intermediate_reg_1[2974]),.o(intermediate_reg_2[1487])); 
xor_module xor_module_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2973]),.i2(intermediate_reg_1[2972]),.o(intermediate_reg_2[1486])); 
xor_module xor_module_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2971]),.i2(intermediate_reg_1[2970]),.o(intermediate_reg_2[1485])); 
mux_module mux_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2969]),.i2(intermediate_reg_1[2968]),.o(intermediate_reg_2[1484]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2967]),.i2(intermediate_reg_1[2966]),.o(intermediate_reg_2[1483])); 
mux_module mux_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2965]),.i2(intermediate_reg_1[2964]),.o(intermediate_reg_2[1482]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2963]),.i2(intermediate_reg_1[2962]),.o(intermediate_reg_2[1481])); 
xor_module xor_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2961]),.i2(intermediate_reg_1[2960]),.o(intermediate_reg_2[1480])); 
xor_module xor_module_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2959]),.i2(intermediate_reg_1[2958]),.o(intermediate_reg_2[1479])); 
xor_module xor_module_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2957]),.i2(intermediate_reg_1[2956]),.o(intermediate_reg_2[1478])); 
xor_module xor_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2955]),.i2(intermediate_reg_1[2954]),.o(intermediate_reg_2[1477])); 
mux_module mux_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2953]),.i2(intermediate_reg_1[2952]),.o(intermediate_reg_2[1476]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2951]),.i2(intermediate_reg_1[2950]),.o(intermediate_reg_2[1475]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2949]),.i2(intermediate_reg_1[2948]),.o(intermediate_reg_2[1474]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2947]),.i2(intermediate_reg_1[2946]),.o(intermediate_reg_2[1473]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2945]),.i2(intermediate_reg_1[2944]),.o(intermediate_reg_2[1472]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2943]),.i2(intermediate_reg_1[2942]),.o(intermediate_reg_2[1471])); 
xor_module xor_module_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2941]),.i2(intermediate_reg_1[2940]),.o(intermediate_reg_2[1470])); 
mux_module mux_module_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2939]),.i2(intermediate_reg_1[2938]),.o(intermediate_reg_2[1469]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2937]),.i2(intermediate_reg_1[2936]),.o(intermediate_reg_2[1468])); 
mux_module mux_module_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2935]),.i2(intermediate_reg_1[2934]),.o(intermediate_reg_2[1467]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2933]),.i2(intermediate_reg_1[2932]),.o(intermediate_reg_2[1466]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2931]),.i2(intermediate_reg_1[2930]),.o(intermediate_reg_2[1465]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2929]),.i2(intermediate_reg_1[2928]),.o(intermediate_reg_2[1464]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2927]),.i2(intermediate_reg_1[2926]),.o(intermediate_reg_2[1463])); 
mux_module mux_module_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2925]),.i2(intermediate_reg_1[2924]),.o(intermediate_reg_2[1462]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2923]),.i2(intermediate_reg_1[2922]),.o(intermediate_reg_2[1461]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2921]),.i2(intermediate_reg_1[2920]),.o(intermediate_reg_2[1460]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2919]),.i2(intermediate_reg_1[2918]),.o(intermediate_reg_2[1459]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2917]),.i2(intermediate_reg_1[2916]),.o(intermediate_reg_2[1458]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2915]),.i2(intermediate_reg_1[2914]),.o(intermediate_reg_2[1457]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2913]),.i2(intermediate_reg_1[2912]),.o(intermediate_reg_2[1456]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2911]),.i2(intermediate_reg_1[2910]),.o(intermediate_reg_2[1455]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2909]),.i2(intermediate_reg_1[2908]),.o(intermediate_reg_2[1454]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2907]),.i2(intermediate_reg_1[2906]),.o(intermediate_reg_2[1453])); 
xor_module xor_module_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2905]),.i2(intermediate_reg_1[2904]),.o(intermediate_reg_2[1452])); 
mux_module mux_module_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2903]),.i2(intermediate_reg_1[2902]),.o(intermediate_reg_2[1451]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2901]),.i2(intermediate_reg_1[2900]),.o(intermediate_reg_2[1450])); 
mux_module mux_module_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2899]),.i2(intermediate_reg_1[2898]),.o(intermediate_reg_2[1449]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2897]),.i2(intermediate_reg_1[2896]),.o(intermediate_reg_2[1448]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2895]),.i2(intermediate_reg_1[2894]),.o(intermediate_reg_2[1447])); 
xor_module xor_module_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2893]),.i2(intermediate_reg_1[2892]),.o(intermediate_reg_2[1446])); 
xor_module xor_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2891]),.i2(intermediate_reg_1[2890]),.o(intermediate_reg_2[1445])); 
mux_module mux_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2889]),.i2(intermediate_reg_1[2888]),.o(intermediate_reg_2[1444]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2887]),.i2(intermediate_reg_1[2886]),.o(intermediate_reg_2[1443])); 
xor_module xor_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2885]),.i2(intermediate_reg_1[2884]),.o(intermediate_reg_2[1442])); 
xor_module xor_module_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2883]),.i2(intermediate_reg_1[2882]),.o(intermediate_reg_2[1441])); 
xor_module xor_module_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2881]),.i2(intermediate_reg_1[2880]),.o(intermediate_reg_2[1440])); 
xor_module xor_module_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2879]),.i2(intermediate_reg_1[2878]),.o(intermediate_reg_2[1439])); 
xor_module xor_module_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2877]),.i2(intermediate_reg_1[2876]),.o(intermediate_reg_2[1438])); 
mux_module mux_module_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2875]),.i2(intermediate_reg_1[2874]),.o(intermediate_reg_2[1437]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2873]),.i2(intermediate_reg_1[2872]),.o(intermediate_reg_2[1436])); 
mux_module mux_module_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2871]),.i2(intermediate_reg_1[2870]),.o(intermediate_reg_2[1435]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2869]),.i2(intermediate_reg_1[2868]),.o(intermediate_reg_2[1434]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2867]),.i2(intermediate_reg_1[2866]),.o(intermediate_reg_2[1433])); 
mux_module mux_module_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2865]),.i2(intermediate_reg_1[2864]),.o(intermediate_reg_2[1432]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2863]),.i2(intermediate_reg_1[2862]),.o(intermediate_reg_2[1431]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2861]),.i2(intermediate_reg_1[2860]),.o(intermediate_reg_2[1430]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2859]),.i2(intermediate_reg_1[2858]),.o(intermediate_reg_2[1429])); 
mux_module mux_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2857]),.i2(intermediate_reg_1[2856]),.o(intermediate_reg_2[1428]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2855]),.i2(intermediate_reg_1[2854]),.o(intermediate_reg_2[1427])); 
mux_module mux_module_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2853]),.i2(intermediate_reg_1[2852]),.o(intermediate_reg_2[1426]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2851]),.i2(intermediate_reg_1[2850]),.o(intermediate_reg_2[1425]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2849]),.i2(intermediate_reg_1[2848]),.o(intermediate_reg_2[1424]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2847]),.i2(intermediate_reg_1[2846]),.o(intermediate_reg_2[1423]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2845]),.i2(intermediate_reg_1[2844]),.o(intermediate_reg_2[1422]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2843]),.i2(intermediate_reg_1[2842]),.o(intermediate_reg_2[1421])); 
mux_module mux_module_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2841]),.i2(intermediate_reg_1[2840]),.o(intermediate_reg_2[1420]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2839]),.i2(intermediate_reg_1[2838]),.o(intermediate_reg_2[1419]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2837]),.i2(intermediate_reg_1[2836]),.o(intermediate_reg_2[1418])); 
mux_module mux_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2835]),.i2(intermediate_reg_1[2834]),.o(intermediate_reg_2[1417]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2833]),.i2(intermediate_reg_1[2832]),.o(intermediate_reg_2[1416]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2831]),.i2(intermediate_reg_1[2830]),.o(intermediate_reg_2[1415])); 
mux_module mux_module_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2829]),.i2(intermediate_reg_1[2828]),.o(intermediate_reg_2[1414]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2827]),.i2(intermediate_reg_1[2826]),.o(intermediate_reg_2[1413])); 
mux_module mux_module_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2825]),.i2(intermediate_reg_1[2824]),.o(intermediate_reg_2[1412]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2823]),.i2(intermediate_reg_1[2822]),.o(intermediate_reg_2[1411]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2821]),.i2(intermediate_reg_1[2820]),.o(intermediate_reg_2[1410]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2819]),.i2(intermediate_reg_1[2818]),.o(intermediate_reg_2[1409]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2817]),.i2(intermediate_reg_1[2816]),.o(intermediate_reg_2[1408]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2815]),.i2(intermediate_reg_1[2814]),.o(intermediate_reg_2[1407]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2813]),.i2(intermediate_reg_1[2812]),.o(intermediate_reg_2[1406]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2811]),.i2(intermediate_reg_1[2810]),.o(intermediate_reg_2[1405])); 
xor_module xor_module_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2809]),.i2(intermediate_reg_1[2808]),.o(intermediate_reg_2[1404])); 
mux_module mux_module_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2807]),.i2(intermediate_reg_1[2806]),.o(intermediate_reg_2[1403]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2805]),.i2(intermediate_reg_1[2804]),.o(intermediate_reg_2[1402])); 
mux_module mux_module_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2803]),.i2(intermediate_reg_1[2802]),.o(intermediate_reg_2[1401]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2801]),.i2(intermediate_reg_1[2800]),.o(intermediate_reg_2[1400])); 
xor_module xor_module_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2799]),.i2(intermediate_reg_1[2798]),.o(intermediate_reg_2[1399])); 
mux_module mux_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2797]),.i2(intermediate_reg_1[2796]),.o(intermediate_reg_2[1398]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2795]),.i2(intermediate_reg_1[2794]),.o(intermediate_reg_2[1397])); 
xor_module xor_module_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2793]),.i2(intermediate_reg_1[2792]),.o(intermediate_reg_2[1396])); 
mux_module mux_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2791]),.i2(intermediate_reg_1[2790]),.o(intermediate_reg_2[1395]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2789]),.i2(intermediate_reg_1[2788]),.o(intermediate_reg_2[1394]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2787]),.i2(intermediate_reg_1[2786]),.o(intermediate_reg_2[1393]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2785]),.i2(intermediate_reg_1[2784]),.o(intermediate_reg_2[1392]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2783]),.i2(intermediate_reg_1[2782]),.o(intermediate_reg_2[1391])); 
xor_module xor_module_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2781]),.i2(intermediate_reg_1[2780]),.o(intermediate_reg_2[1390])); 
xor_module xor_module_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2779]),.i2(intermediate_reg_1[2778]),.o(intermediate_reg_2[1389])); 
mux_module mux_module_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2777]),.i2(intermediate_reg_1[2776]),.o(intermediate_reg_2[1388]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2775]),.i2(intermediate_reg_1[2774]),.o(intermediate_reg_2[1387])); 
xor_module xor_module_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2773]),.i2(intermediate_reg_1[2772]),.o(intermediate_reg_2[1386])); 
xor_module xor_module_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2771]),.i2(intermediate_reg_1[2770]),.o(intermediate_reg_2[1385])); 
mux_module mux_module_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2769]),.i2(intermediate_reg_1[2768]),.o(intermediate_reg_2[1384]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2767]),.i2(intermediate_reg_1[2766]),.o(intermediate_reg_2[1383])); 
mux_module mux_module_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2765]),.i2(intermediate_reg_1[2764]),.o(intermediate_reg_2[1382]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2763]),.i2(intermediate_reg_1[2762]),.o(intermediate_reg_2[1381])); 
xor_module xor_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2761]),.i2(intermediate_reg_1[2760]),.o(intermediate_reg_2[1380])); 
mux_module mux_module_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2759]),.i2(intermediate_reg_1[2758]),.o(intermediate_reg_2[1379]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2757]),.i2(intermediate_reg_1[2756]),.o(intermediate_reg_2[1378]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2755]),.i2(intermediate_reg_1[2754]),.o(intermediate_reg_2[1377]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2753]),.i2(intermediate_reg_1[2752]),.o(intermediate_reg_2[1376])); 
mux_module mux_module_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2751]),.i2(intermediate_reg_1[2750]),.o(intermediate_reg_2[1375]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2749]),.i2(intermediate_reg_1[2748]),.o(intermediate_reg_2[1374])); 
xor_module xor_module_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2747]),.i2(intermediate_reg_1[2746]),.o(intermediate_reg_2[1373])); 
mux_module mux_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2745]),.i2(intermediate_reg_1[2744]),.o(intermediate_reg_2[1372]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2743]),.i2(intermediate_reg_1[2742]),.o(intermediate_reg_2[1371])); 
xor_module xor_module_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2741]),.i2(intermediate_reg_1[2740]),.o(intermediate_reg_2[1370])); 
mux_module mux_module_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2739]),.i2(intermediate_reg_1[2738]),.o(intermediate_reg_2[1369]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2737]),.i2(intermediate_reg_1[2736]),.o(intermediate_reg_2[1368]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2735]),.i2(intermediate_reg_1[2734]),.o(intermediate_reg_2[1367]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2733]),.i2(intermediate_reg_1[2732]),.o(intermediate_reg_2[1366]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2731]),.i2(intermediate_reg_1[2730]),.o(intermediate_reg_2[1365]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2729]),.i2(intermediate_reg_1[2728]),.o(intermediate_reg_2[1364])); 
mux_module mux_module_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2727]),.i2(intermediate_reg_1[2726]),.o(intermediate_reg_2[1363]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2725]),.i2(intermediate_reg_1[2724]),.o(intermediate_reg_2[1362])); 
xor_module xor_module_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2723]),.i2(intermediate_reg_1[2722]),.o(intermediate_reg_2[1361])); 
mux_module mux_module_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2721]),.i2(intermediate_reg_1[2720]),.o(intermediate_reg_2[1360]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2719]),.i2(intermediate_reg_1[2718]),.o(intermediate_reg_2[1359])); 
xor_module xor_module_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2717]),.i2(intermediate_reg_1[2716]),.o(intermediate_reg_2[1358])); 
xor_module xor_module_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2715]),.i2(intermediate_reg_1[2714]),.o(intermediate_reg_2[1357])); 
mux_module mux_module_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2713]),.i2(intermediate_reg_1[2712]),.o(intermediate_reg_2[1356]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2711]),.i2(intermediate_reg_1[2710]),.o(intermediate_reg_2[1355]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2709]),.i2(intermediate_reg_1[2708]),.o(intermediate_reg_2[1354]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2707]),.i2(intermediate_reg_1[2706]),.o(intermediate_reg_2[1353])); 
xor_module xor_module_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2705]),.i2(intermediate_reg_1[2704]),.o(intermediate_reg_2[1352])); 
mux_module mux_module_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2703]),.i2(intermediate_reg_1[2702]),.o(intermediate_reg_2[1351]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2701]),.i2(intermediate_reg_1[2700]),.o(intermediate_reg_2[1350])); 
xor_module xor_module_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2699]),.i2(intermediate_reg_1[2698]),.o(intermediate_reg_2[1349])); 
mux_module mux_module_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2697]),.i2(intermediate_reg_1[2696]),.o(intermediate_reg_2[1348]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2695]),.i2(intermediate_reg_1[2694]),.o(intermediate_reg_2[1347]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2693]),.i2(intermediate_reg_1[2692]),.o(intermediate_reg_2[1346]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2691]),.i2(intermediate_reg_1[2690]),.o(intermediate_reg_2[1345])); 
xor_module xor_module_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2689]),.i2(intermediate_reg_1[2688]),.o(intermediate_reg_2[1344])); 
mux_module mux_module_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2687]),.i2(intermediate_reg_1[2686]),.o(intermediate_reg_2[1343]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2685]),.i2(intermediate_reg_1[2684]),.o(intermediate_reg_2[1342])); 
xor_module xor_module_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2683]),.i2(intermediate_reg_1[2682]),.o(intermediate_reg_2[1341])); 
xor_module xor_module_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2681]),.i2(intermediate_reg_1[2680]),.o(intermediate_reg_2[1340])); 
mux_module mux_module_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2679]),.i2(intermediate_reg_1[2678]),.o(intermediate_reg_2[1339]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2677]),.i2(intermediate_reg_1[2676]),.o(intermediate_reg_2[1338])); 
xor_module xor_module_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2675]),.i2(intermediate_reg_1[2674]),.o(intermediate_reg_2[1337])); 
xor_module xor_module_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2673]),.i2(intermediate_reg_1[2672]),.o(intermediate_reg_2[1336])); 
mux_module mux_module_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2671]),.i2(intermediate_reg_1[2670]),.o(intermediate_reg_2[1335]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2669]),.i2(intermediate_reg_1[2668]),.o(intermediate_reg_2[1334]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2667]),.i2(intermediate_reg_1[2666]),.o(intermediate_reg_2[1333])); 
mux_module mux_module_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2665]),.i2(intermediate_reg_1[2664]),.o(intermediate_reg_2[1332]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2663]),.i2(intermediate_reg_1[2662]),.o(intermediate_reg_2[1331])); 
mux_module mux_module_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2661]),.i2(intermediate_reg_1[2660]),.o(intermediate_reg_2[1330]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2659]),.i2(intermediate_reg_1[2658]),.o(intermediate_reg_2[1329]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2657]),.i2(intermediate_reg_1[2656]),.o(intermediate_reg_2[1328]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2655]),.i2(intermediate_reg_1[2654]),.o(intermediate_reg_2[1327]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2653]),.i2(intermediate_reg_1[2652]),.o(intermediate_reg_2[1326])); 
xor_module xor_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2651]),.i2(intermediate_reg_1[2650]),.o(intermediate_reg_2[1325])); 
xor_module xor_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2649]),.i2(intermediate_reg_1[2648]),.o(intermediate_reg_2[1324])); 
xor_module xor_module_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2647]),.i2(intermediate_reg_1[2646]),.o(intermediate_reg_2[1323])); 
mux_module mux_module_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2645]),.i2(intermediate_reg_1[2644]),.o(intermediate_reg_2[1322]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2643]),.i2(intermediate_reg_1[2642]),.o(intermediate_reg_2[1321]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2641]),.i2(intermediate_reg_1[2640]),.o(intermediate_reg_2[1320]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2639]),.i2(intermediate_reg_1[2638]),.o(intermediate_reg_2[1319])); 
xor_module xor_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2637]),.i2(intermediate_reg_1[2636]),.o(intermediate_reg_2[1318])); 
mux_module mux_module_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2635]),.i2(intermediate_reg_1[2634]),.o(intermediate_reg_2[1317]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2633]),.i2(intermediate_reg_1[2632]),.o(intermediate_reg_2[1316]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2631]),.i2(intermediate_reg_1[2630]),.o(intermediate_reg_2[1315]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2629]),.i2(intermediate_reg_1[2628]),.o(intermediate_reg_2[1314])); 
mux_module mux_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2627]),.i2(intermediate_reg_1[2626]),.o(intermediate_reg_2[1313]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2625]),.i2(intermediate_reg_1[2624]),.o(intermediate_reg_2[1312]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2623]),.i2(intermediate_reg_1[2622]),.o(intermediate_reg_2[1311]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2621]),.i2(intermediate_reg_1[2620]),.o(intermediate_reg_2[1310])); 
mux_module mux_module_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2619]),.i2(intermediate_reg_1[2618]),.o(intermediate_reg_2[1309]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2617]),.i2(intermediate_reg_1[2616]),.o(intermediate_reg_2[1308]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2615]),.i2(intermediate_reg_1[2614]),.o(intermediate_reg_2[1307])); 
mux_module mux_module_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2613]),.i2(intermediate_reg_1[2612]),.o(intermediate_reg_2[1306]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2611]),.i2(intermediate_reg_1[2610]),.o(intermediate_reg_2[1305]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2609]),.i2(intermediate_reg_1[2608]),.o(intermediate_reg_2[1304])); 
mux_module mux_module_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2607]),.i2(intermediate_reg_1[2606]),.o(intermediate_reg_2[1303]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2605]),.i2(intermediate_reg_1[2604]),.o(intermediate_reg_2[1302]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2603]),.i2(intermediate_reg_1[2602]),.o(intermediate_reg_2[1301]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2601]),.i2(intermediate_reg_1[2600]),.o(intermediate_reg_2[1300])); 
xor_module xor_module_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2599]),.i2(intermediate_reg_1[2598]),.o(intermediate_reg_2[1299])); 
mux_module mux_module_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2597]),.i2(intermediate_reg_1[2596]),.o(intermediate_reg_2[1298]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2595]),.i2(intermediate_reg_1[2594]),.o(intermediate_reg_2[1297]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2593]),.i2(intermediate_reg_1[2592]),.o(intermediate_reg_2[1296]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2591]),.i2(intermediate_reg_1[2590]),.o(intermediate_reg_2[1295]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2589]),.i2(intermediate_reg_1[2588]),.o(intermediate_reg_2[1294])); 
mux_module mux_module_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2587]),.i2(intermediate_reg_1[2586]),.o(intermediate_reg_2[1293]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2585]),.i2(intermediate_reg_1[2584]),.o(intermediate_reg_2[1292])); 
xor_module xor_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2583]),.i2(intermediate_reg_1[2582]),.o(intermediate_reg_2[1291])); 
xor_module xor_module_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2581]),.i2(intermediate_reg_1[2580]),.o(intermediate_reg_2[1290])); 
xor_module xor_module_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2579]),.i2(intermediate_reg_1[2578]),.o(intermediate_reg_2[1289])); 
xor_module xor_module_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2577]),.i2(intermediate_reg_1[2576]),.o(intermediate_reg_2[1288])); 
xor_module xor_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2575]),.i2(intermediate_reg_1[2574]),.o(intermediate_reg_2[1287])); 
xor_module xor_module_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2573]),.i2(intermediate_reg_1[2572]),.o(intermediate_reg_2[1286])); 
xor_module xor_module_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2571]),.i2(intermediate_reg_1[2570]),.o(intermediate_reg_2[1285])); 
xor_module xor_module_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2569]),.i2(intermediate_reg_1[2568]),.o(intermediate_reg_2[1284])); 
mux_module mux_module_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2567]),.i2(intermediate_reg_1[2566]),.o(intermediate_reg_2[1283]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2565]),.i2(intermediate_reg_1[2564]),.o(intermediate_reg_2[1282]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2563]),.i2(intermediate_reg_1[2562]),.o(intermediate_reg_2[1281]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2561]),.i2(intermediate_reg_1[2560]),.o(intermediate_reg_2[1280])); 
mux_module mux_module_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2559]),.i2(intermediate_reg_1[2558]),.o(intermediate_reg_2[1279]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2557]),.i2(intermediate_reg_1[2556]),.o(intermediate_reg_2[1278])); 
mux_module mux_module_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2555]),.i2(intermediate_reg_1[2554]),.o(intermediate_reg_2[1277]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2553]),.i2(intermediate_reg_1[2552]),.o(intermediate_reg_2[1276]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2551]),.i2(intermediate_reg_1[2550]),.o(intermediate_reg_2[1275]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2549]),.i2(intermediate_reg_1[2548]),.o(intermediate_reg_2[1274]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2547]),.i2(intermediate_reg_1[2546]),.o(intermediate_reg_2[1273]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2545]),.i2(intermediate_reg_1[2544]),.o(intermediate_reg_2[1272]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2543]),.i2(intermediate_reg_1[2542]),.o(intermediate_reg_2[1271]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2541]),.i2(intermediate_reg_1[2540]),.o(intermediate_reg_2[1270])); 
xor_module xor_module_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2539]),.i2(intermediate_reg_1[2538]),.o(intermediate_reg_2[1269])); 
xor_module xor_module_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2537]),.i2(intermediate_reg_1[2536]),.o(intermediate_reg_2[1268])); 
xor_module xor_module_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2535]),.i2(intermediate_reg_1[2534]),.o(intermediate_reg_2[1267])); 
mux_module mux_module_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2533]),.i2(intermediate_reg_1[2532]),.o(intermediate_reg_2[1266]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2531]),.i2(intermediate_reg_1[2530]),.o(intermediate_reg_2[1265])); 
mux_module mux_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2529]),.i2(intermediate_reg_1[2528]),.o(intermediate_reg_2[1264]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2527]),.i2(intermediate_reg_1[2526]),.o(intermediate_reg_2[1263])); 
xor_module xor_module_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2525]),.i2(intermediate_reg_1[2524]),.o(intermediate_reg_2[1262])); 
mux_module mux_module_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2523]),.i2(intermediate_reg_1[2522]),.o(intermediate_reg_2[1261]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2521]),.i2(intermediate_reg_1[2520]),.o(intermediate_reg_2[1260])); 
mux_module mux_module_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2519]),.i2(intermediate_reg_1[2518]),.o(intermediate_reg_2[1259]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2517]),.i2(intermediate_reg_1[2516]),.o(intermediate_reg_2[1258])); 
xor_module xor_module_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2515]),.i2(intermediate_reg_1[2514]),.o(intermediate_reg_2[1257])); 
mux_module mux_module_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2513]),.i2(intermediate_reg_1[2512]),.o(intermediate_reg_2[1256]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2511]),.i2(intermediate_reg_1[2510]),.o(intermediate_reg_2[1255]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2509]),.i2(intermediate_reg_1[2508]),.o(intermediate_reg_2[1254])); 
xor_module xor_module_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2507]),.i2(intermediate_reg_1[2506]),.o(intermediate_reg_2[1253])); 
xor_module xor_module_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2505]),.i2(intermediate_reg_1[2504]),.o(intermediate_reg_2[1252])); 
xor_module xor_module_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2503]),.i2(intermediate_reg_1[2502]),.o(intermediate_reg_2[1251])); 
xor_module xor_module_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2501]),.i2(intermediate_reg_1[2500]),.o(intermediate_reg_2[1250])); 
mux_module mux_module_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2499]),.i2(intermediate_reg_1[2498]),.o(intermediate_reg_2[1249]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2497]),.i2(intermediate_reg_1[2496]),.o(intermediate_reg_2[1248]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2495]),.i2(intermediate_reg_1[2494]),.o(intermediate_reg_2[1247]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2493]),.i2(intermediate_reg_1[2492]),.o(intermediate_reg_2[1246])); 
xor_module xor_module_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2491]),.i2(intermediate_reg_1[2490]),.o(intermediate_reg_2[1245])); 
mux_module mux_module_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2489]),.i2(intermediate_reg_1[2488]),.o(intermediate_reg_2[1244]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2487]),.i2(intermediate_reg_1[2486]),.o(intermediate_reg_2[1243])); 
mux_module mux_module_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2485]),.i2(intermediate_reg_1[2484]),.o(intermediate_reg_2[1242]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2483]),.i2(intermediate_reg_1[2482]),.o(intermediate_reg_2[1241]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2481]),.i2(intermediate_reg_1[2480]),.o(intermediate_reg_2[1240])); 
mux_module mux_module_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2479]),.i2(intermediate_reg_1[2478]),.o(intermediate_reg_2[1239]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2477]),.i2(intermediate_reg_1[2476]),.o(intermediate_reg_2[1238])); 
xor_module xor_module_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2475]),.i2(intermediate_reg_1[2474]),.o(intermediate_reg_2[1237])); 
xor_module xor_module_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2473]),.i2(intermediate_reg_1[2472]),.o(intermediate_reg_2[1236])); 
mux_module mux_module_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2471]),.i2(intermediate_reg_1[2470]),.o(intermediate_reg_2[1235]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2469]),.i2(intermediate_reg_1[2468]),.o(intermediate_reg_2[1234]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2467]),.i2(intermediate_reg_1[2466]),.o(intermediate_reg_2[1233]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2465]),.i2(intermediate_reg_1[2464]),.o(intermediate_reg_2[1232]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2463]),.i2(intermediate_reg_1[2462]),.o(intermediate_reg_2[1231]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2461]),.i2(intermediate_reg_1[2460]),.o(intermediate_reg_2[1230])); 
mux_module mux_module_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2459]),.i2(intermediate_reg_1[2458]),.o(intermediate_reg_2[1229]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2457]),.i2(intermediate_reg_1[2456]),.o(intermediate_reg_2[1228])); 
xor_module xor_module_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2455]),.i2(intermediate_reg_1[2454]),.o(intermediate_reg_2[1227])); 
xor_module xor_module_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2453]),.i2(intermediate_reg_1[2452]),.o(intermediate_reg_2[1226])); 
mux_module mux_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2451]),.i2(intermediate_reg_1[2450]),.o(intermediate_reg_2[1225]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2449]),.i2(intermediate_reg_1[2448]),.o(intermediate_reg_2[1224])); 
xor_module xor_module_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2447]),.i2(intermediate_reg_1[2446]),.o(intermediate_reg_2[1223])); 
xor_module xor_module_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2445]),.i2(intermediate_reg_1[2444]),.o(intermediate_reg_2[1222])); 
mux_module mux_module_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2443]),.i2(intermediate_reg_1[2442]),.o(intermediate_reg_2[1221]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2441]),.i2(intermediate_reg_1[2440]),.o(intermediate_reg_2[1220])); 
xor_module xor_module_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2439]),.i2(intermediate_reg_1[2438]),.o(intermediate_reg_2[1219])); 
xor_module xor_module_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2437]),.i2(intermediate_reg_1[2436]),.o(intermediate_reg_2[1218])); 
xor_module xor_module_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2435]),.i2(intermediate_reg_1[2434]),.o(intermediate_reg_2[1217])); 
xor_module xor_module_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2433]),.i2(intermediate_reg_1[2432]),.o(intermediate_reg_2[1216])); 
xor_module xor_module_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2431]),.i2(intermediate_reg_1[2430]),.o(intermediate_reg_2[1215])); 
mux_module mux_module_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2429]),.i2(intermediate_reg_1[2428]),.o(intermediate_reg_2[1214]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2427]),.i2(intermediate_reg_1[2426]),.o(intermediate_reg_2[1213]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2425]),.i2(intermediate_reg_1[2424]),.o(intermediate_reg_2[1212]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2423]),.i2(intermediate_reg_1[2422]),.o(intermediate_reg_2[1211]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2421]),.i2(intermediate_reg_1[2420]),.o(intermediate_reg_2[1210]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2419]),.i2(intermediate_reg_1[2418]),.o(intermediate_reg_2[1209]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2417]),.i2(intermediate_reg_1[2416]),.o(intermediate_reg_2[1208]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2415]),.i2(intermediate_reg_1[2414]),.o(intermediate_reg_2[1207])); 
xor_module xor_module_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2413]),.i2(intermediate_reg_1[2412]),.o(intermediate_reg_2[1206])); 
mux_module mux_module_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2411]),.i2(intermediate_reg_1[2410]),.o(intermediate_reg_2[1205]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2409]),.i2(intermediate_reg_1[2408]),.o(intermediate_reg_2[1204])); 
xor_module xor_module_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2407]),.i2(intermediate_reg_1[2406]),.o(intermediate_reg_2[1203])); 
mux_module mux_module_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2405]),.i2(intermediate_reg_1[2404]),.o(intermediate_reg_2[1202]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2403]),.i2(intermediate_reg_1[2402]),.o(intermediate_reg_2[1201])); 
xor_module xor_module_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2401]),.i2(intermediate_reg_1[2400]),.o(intermediate_reg_2[1200])); 
xor_module xor_module_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2399]),.i2(intermediate_reg_1[2398]),.o(intermediate_reg_2[1199])); 
xor_module xor_module_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2397]),.i2(intermediate_reg_1[2396]),.o(intermediate_reg_2[1198])); 
xor_module xor_module_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2395]),.i2(intermediate_reg_1[2394]),.o(intermediate_reg_2[1197])); 
xor_module xor_module_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2393]),.i2(intermediate_reg_1[2392]),.o(intermediate_reg_2[1196])); 
xor_module xor_module_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2391]),.i2(intermediate_reg_1[2390]),.o(intermediate_reg_2[1195])); 
xor_module xor_module_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2389]),.i2(intermediate_reg_1[2388]),.o(intermediate_reg_2[1194])); 
mux_module mux_module_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2387]),.i2(intermediate_reg_1[2386]),.o(intermediate_reg_2[1193]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2385]),.i2(intermediate_reg_1[2384]),.o(intermediate_reg_2[1192]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2383]),.i2(intermediate_reg_1[2382]),.o(intermediate_reg_2[1191])); 
mux_module mux_module_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2381]),.i2(intermediate_reg_1[2380]),.o(intermediate_reg_2[1190]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2379]),.i2(intermediate_reg_1[2378]),.o(intermediate_reg_2[1189])); 
mux_module mux_module_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2377]),.i2(intermediate_reg_1[2376]),.o(intermediate_reg_2[1188]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2375]),.i2(intermediate_reg_1[2374]),.o(intermediate_reg_2[1187])); 
mux_module mux_module_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2373]),.i2(intermediate_reg_1[2372]),.o(intermediate_reg_2[1186]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2371]),.i2(intermediate_reg_1[2370]),.o(intermediate_reg_2[1185])); 
mux_module mux_module_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2369]),.i2(intermediate_reg_1[2368]),.o(intermediate_reg_2[1184]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2367]),.i2(intermediate_reg_1[2366]),.o(intermediate_reg_2[1183]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2365]),.i2(intermediate_reg_1[2364]),.o(intermediate_reg_2[1182])); 
mux_module mux_module_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2363]),.i2(intermediate_reg_1[2362]),.o(intermediate_reg_2[1181]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2361]),.i2(intermediate_reg_1[2360]),.o(intermediate_reg_2[1180])); 
mux_module mux_module_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2359]),.i2(intermediate_reg_1[2358]),.o(intermediate_reg_2[1179]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2357]),.i2(intermediate_reg_1[2356]),.o(intermediate_reg_2[1178]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2355]),.i2(intermediate_reg_1[2354]),.o(intermediate_reg_2[1177])); 
mux_module mux_module_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2353]),.i2(intermediate_reg_1[2352]),.o(intermediate_reg_2[1176]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2351]),.i2(intermediate_reg_1[2350]),.o(intermediate_reg_2[1175]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2349]),.i2(intermediate_reg_1[2348]),.o(intermediate_reg_2[1174])); 
mux_module mux_module_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2347]),.i2(intermediate_reg_1[2346]),.o(intermediate_reg_2[1173]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2345]),.i2(intermediate_reg_1[2344]),.o(intermediate_reg_2[1172]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2343]),.i2(intermediate_reg_1[2342]),.o(intermediate_reg_2[1171])); 
mux_module mux_module_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2341]),.i2(intermediate_reg_1[2340]),.o(intermediate_reg_2[1170]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2339]),.i2(intermediate_reg_1[2338]),.o(intermediate_reg_2[1169])); 
xor_module xor_module_inst_2_480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2337]),.i2(intermediate_reg_1[2336]),.o(intermediate_reg_2[1168])); 
xor_module xor_module_inst_2_481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2335]),.i2(intermediate_reg_1[2334]),.o(intermediate_reg_2[1167])); 
mux_module mux_module_inst_2_482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2333]),.i2(intermediate_reg_1[2332]),.o(intermediate_reg_2[1166]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2331]),.i2(intermediate_reg_1[2330]),.o(intermediate_reg_2[1165]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2329]),.i2(intermediate_reg_1[2328]),.o(intermediate_reg_2[1164])); 
xor_module xor_module_inst_2_485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2327]),.i2(intermediate_reg_1[2326]),.o(intermediate_reg_2[1163])); 
mux_module mux_module_inst_2_486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2325]),.i2(intermediate_reg_1[2324]),.o(intermediate_reg_2[1162]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2323]),.i2(intermediate_reg_1[2322]),.o(intermediate_reg_2[1161])); 
xor_module xor_module_inst_2_488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2321]),.i2(intermediate_reg_1[2320]),.o(intermediate_reg_2[1160])); 
mux_module mux_module_inst_2_489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2319]),.i2(intermediate_reg_1[2318]),.o(intermediate_reg_2[1159]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2317]),.i2(intermediate_reg_1[2316]),.o(intermediate_reg_2[1158])); 
mux_module mux_module_inst_2_491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2315]),.i2(intermediate_reg_1[2314]),.o(intermediate_reg_2[1157]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2313]),.i2(intermediate_reg_1[2312]),.o(intermediate_reg_2[1156]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2311]),.i2(intermediate_reg_1[2310]),.o(intermediate_reg_2[1155]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2309]),.i2(intermediate_reg_1[2308]),.o(intermediate_reg_2[1154])); 
mux_module mux_module_inst_2_495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2307]),.i2(intermediate_reg_1[2306]),.o(intermediate_reg_2[1153]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2305]),.i2(intermediate_reg_1[2304]),.o(intermediate_reg_2[1152]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2303]),.i2(intermediate_reg_1[2302]),.o(intermediate_reg_2[1151])); 
xor_module xor_module_inst_2_498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2301]),.i2(intermediate_reg_1[2300]),.o(intermediate_reg_2[1150])); 
xor_module xor_module_inst_2_499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2299]),.i2(intermediate_reg_1[2298]),.o(intermediate_reg_2[1149])); 
mux_module mux_module_inst_2_500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2297]),.i2(intermediate_reg_1[2296]),.o(intermediate_reg_2[1148]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2295]),.i2(intermediate_reg_1[2294]),.o(intermediate_reg_2[1147])); 
xor_module xor_module_inst_2_502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2293]),.i2(intermediate_reg_1[2292]),.o(intermediate_reg_2[1146])); 
mux_module mux_module_inst_2_503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2291]),.i2(intermediate_reg_1[2290]),.o(intermediate_reg_2[1145]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2289]),.i2(intermediate_reg_1[2288]),.o(intermediate_reg_2[1144]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2287]),.i2(intermediate_reg_1[2286]),.o(intermediate_reg_2[1143])); 
mux_module mux_module_inst_2_506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2285]),.i2(intermediate_reg_1[2284]),.o(intermediate_reg_2[1142]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2283]),.i2(intermediate_reg_1[2282]),.o(intermediate_reg_2[1141]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2281]),.i2(intermediate_reg_1[2280]),.o(intermediate_reg_2[1140]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2279]),.i2(intermediate_reg_1[2278]),.o(intermediate_reg_2[1139])); 
mux_module mux_module_inst_2_510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2277]),.i2(intermediate_reg_1[2276]),.o(intermediate_reg_2[1138]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2275]),.i2(intermediate_reg_1[2274]),.o(intermediate_reg_2[1137]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2273]),.i2(intermediate_reg_1[2272]),.o(intermediate_reg_2[1136]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2271]),.i2(intermediate_reg_1[2270]),.o(intermediate_reg_2[1135])); 
xor_module xor_module_inst_2_514(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2269]),.i2(intermediate_reg_1[2268]),.o(intermediate_reg_2[1134])); 
xor_module xor_module_inst_2_515(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2267]),.i2(intermediate_reg_1[2266]),.o(intermediate_reg_2[1133])); 
mux_module mux_module_inst_2_516(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2265]),.i2(intermediate_reg_1[2264]),.o(intermediate_reg_2[1132]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_517(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2263]),.i2(intermediate_reg_1[2262]),.o(intermediate_reg_2[1131])); 
xor_module xor_module_inst_2_518(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2261]),.i2(intermediate_reg_1[2260]),.o(intermediate_reg_2[1130])); 
xor_module xor_module_inst_2_519(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2259]),.i2(intermediate_reg_1[2258]),.o(intermediate_reg_2[1129])); 
mux_module mux_module_inst_2_520(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2257]),.i2(intermediate_reg_1[2256]),.o(intermediate_reg_2[1128]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_521(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2255]),.i2(intermediate_reg_1[2254]),.o(intermediate_reg_2[1127])); 
xor_module xor_module_inst_2_522(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2253]),.i2(intermediate_reg_1[2252]),.o(intermediate_reg_2[1126])); 
mux_module mux_module_inst_2_523(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2251]),.i2(intermediate_reg_1[2250]),.o(intermediate_reg_2[1125]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_524(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2249]),.i2(intermediate_reg_1[2248]),.o(intermediate_reg_2[1124])); 
mux_module mux_module_inst_2_525(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2247]),.i2(intermediate_reg_1[2246]),.o(intermediate_reg_2[1123]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_526(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2245]),.i2(intermediate_reg_1[2244]),.o(intermediate_reg_2[1122]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_527(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2243]),.i2(intermediate_reg_1[2242]),.o(intermediate_reg_2[1121]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_528(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2241]),.i2(intermediate_reg_1[2240]),.o(intermediate_reg_2[1120])); 
mux_module mux_module_inst_2_529(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2239]),.i2(intermediate_reg_1[2238]),.o(intermediate_reg_2[1119]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_530(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2237]),.i2(intermediate_reg_1[2236]),.o(intermediate_reg_2[1118]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_531(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2235]),.i2(intermediate_reg_1[2234]),.o(intermediate_reg_2[1117])); 
xor_module xor_module_inst_2_532(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2233]),.i2(intermediate_reg_1[2232]),.o(intermediate_reg_2[1116])); 
mux_module mux_module_inst_2_533(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2231]),.i2(intermediate_reg_1[2230]),.o(intermediate_reg_2[1115]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_534(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2229]),.i2(intermediate_reg_1[2228]),.o(intermediate_reg_2[1114]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_535(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2227]),.i2(intermediate_reg_1[2226]),.o(intermediate_reg_2[1113]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_536(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2225]),.i2(intermediate_reg_1[2224]),.o(intermediate_reg_2[1112]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_537(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2223]),.i2(intermediate_reg_1[2222]),.o(intermediate_reg_2[1111]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_538(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2221]),.i2(intermediate_reg_1[2220]),.o(intermediate_reg_2[1110])); 
mux_module mux_module_inst_2_539(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2219]),.i2(intermediate_reg_1[2218]),.o(intermediate_reg_2[1109]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_540(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2217]),.i2(intermediate_reg_1[2216]),.o(intermediate_reg_2[1108])); 
mux_module mux_module_inst_2_541(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2215]),.i2(intermediate_reg_1[2214]),.o(intermediate_reg_2[1107]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_542(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2213]),.i2(intermediate_reg_1[2212]),.o(intermediate_reg_2[1106])); 
xor_module xor_module_inst_2_543(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2211]),.i2(intermediate_reg_1[2210]),.o(intermediate_reg_2[1105])); 
mux_module mux_module_inst_2_544(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2209]),.i2(intermediate_reg_1[2208]),.o(intermediate_reg_2[1104]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_545(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2207]),.i2(intermediate_reg_1[2206]),.o(intermediate_reg_2[1103])); 
xor_module xor_module_inst_2_546(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2205]),.i2(intermediate_reg_1[2204]),.o(intermediate_reg_2[1102])); 
xor_module xor_module_inst_2_547(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2203]),.i2(intermediate_reg_1[2202]),.o(intermediate_reg_2[1101])); 
mux_module mux_module_inst_2_548(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2201]),.i2(intermediate_reg_1[2200]),.o(intermediate_reg_2[1100]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_549(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2199]),.i2(intermediate_reg_1[2198]),.o(intermediate_reg_2[1099]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_550(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2197]),.i2(intermediate_reg_1[2196]),.o(intermediate_reg_2[1098]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_551(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2195]),.i2(intermediate_reg_1[2194]),.o(intermediate_reg_2[1097]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_552(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2193]),.i2(intermediate_reg_1[2192]),.o(intermediate_reg_2[1096]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_553(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2191]),.i2(intermediate_reg_1[2190]),.o(intermediate_reg_2[1095]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_554(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2189]),.i2(intermediate_reg_1[2188]),.o(intermediate_reg_2[1094])); 
mux_module mux_module_inst_2_555(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2187]),.i2(intermediate_reg_1[2186]),.o(intermediate_reg_2[1093]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_556(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2185]),.i2(intermediate_reg_1[2184]),.o(intermediate_reg_2[1092])); 
mux_module mux_module_inst_2_557(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2183]),.i2(intermediate_reg_1[2182]),.o(intermediate_reg_2[1091]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_558(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2181]),.i2(intermediate_reg_1[2180]),.o(intermediate_reg_2[1090])); 
xor_module xor_module_inst_2_559(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2179]),.i2(intermediate_reg_1[2178]),.o(intermediate_reg_2[1089])); 
xor_module xor_module_inst_2_560(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2177]),.i2(intermediate_reg_1[2176]),.o(intermediate_reg_2[1088])); 
mux_module mux_module_inst_2_561(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2175]),.i2(intermediate_reg_1[2174]),.o(intermediate_reg_2[1087]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_562(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2173]),.i2(intermediate_reg_1[2172]),.o(intermediate_reg_2[1086]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_563(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2171]),.i2(intermediate_reg_1[2170]),.o(intermediate_reg_2[1085])); 
xor_module xor_module_inst_2_564(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2169]),.i2(intermediate_reg_1[2168]),.o(intermediate_reg_2[1084])); 
mux_module mux_module_inst_2_565(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2167]),.i2(intermediate_reg_1[2166]),.o(intermediate_reg_2[1083]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_566(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2165]),.i2(intermediate_reg_1[2164]),.o(intermediate_reg_2[1082])); 
mux_module mux_module_inst_2_567(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2163]),.i2(intermediate_reg_1[2162]),.o(intermediate_reg_2[1081]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_568(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2161]),.i2(intermediate_reg_1[2160]),.o(intermediate_reg_2[1080]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_569(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2159]),.i2(intermediate_reg_1[2158]),.o(intermediate_reg_2[1079]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_570(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2157]),.i2(intermediate_reg_1[2156]),.o(intermediate_reg_2[1078])); 
mux_module mux_module_inst_2_571(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2155]),.i2(intermediate_reg_1[2154]),.o(intermediate_reg_2[1077]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_572(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2153]),.i2(intermediate_reg_1[2152]),.o(intermediate_reg_2[1076]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_573(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2151]),.i2(intermediate_reg_1[2150]),.o(intermediate_reg_2[1075]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_574(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2149]),.i2(intermediate_reg_1[2148]),.o(intermediate_reg_2[1074])); 
mux_module mux_module_inst_2_575(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2147]),.i2(intermediate_reg_1[2146]),.o(intermediate_reg_2[1073]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_576(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2145]),.i2(intermediate_reg_1[2144]),.o(intermediate_reg_2[1072]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_577(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2143]),.i2(intermediate_reg_1[2142]),.o(intermediate_reg_2[1071]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_578(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2141]),.i2(intermediate_reg_1[2140]),.o(intermediate_reg_2[1070])); 
mux_module mux_module_inst_2_579(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2139]),.i2(intermediate_reg_1[2138]),.o(intermediate_reg_2[1069]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_580(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2137]),.i2(intermediate_reg_1[2136]),.o(intermediate_reg_2[1068]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_581(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2135]),.i2(intermediate_reg_1[2134]),.o(intermediate_reg_2[1067]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_582(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2133]),.i2(intermediate_reg_1[2132]),.o(intermediate_reg_2[1066]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_583(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2131]),.i2(intermediate_reg_1[2130]),.o(intermediate_reg_2[1065]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_584(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2129]),.i2(intermediate_reg_1[2128]),.o(intermediate_reg_2[1064])); 
mux_module mux_module_inst_2_585(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2127]),.i2(intermediate_reg_1[2126]),.o(intermediate_reg_2[1063]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_586(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2125]),.i2(intermediate_reg_1[2124]),.o(intermediate_reg_2[1062]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_587(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2123]),.i2(intermediate_reg_1[2122]),.o(intermediate_reg_2[1061])); 
mux_module mux_module_inst_2_588(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2121]),.i2(intermediate_reg_1[2120]),.o(intermediate_reg_2[1060]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_589(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2119]),.i2(intermediate_reg_1[2118]),.o(intermediate_reg_2[1059])); 
xor_module xor_module_inst_2_590(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2117]),.i2(intermediate_reg_1[2116]),.o(intermediate_reg_2[1058])); 
xor_module xor_module_inst_2_591(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2115]),.i2(intermediate_reg_1[2114]),.o(intermediate_reg_2[1057])); 
xor_module xor_module_inst_2_592(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2113]),.i2(intermediate_reg_1[2112]),.o(intermediate_reg_2[1056])); 
xor_module xor_module_inst_2_593(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2111]),.i2(intermediate_reg_1[2110]),.o(intermediate_reg_2[1055])); 
xor_module xor_module_inst_2_594(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2109]),.i2(intermediate_reg_1[2108]),.o(intermediate_reg_2[1054])); 
xor_module xor_module_inst_2_595(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2107]),.i2(intermediate_reg_1[2106]),.o(intermediate_reg_2[1053])); 
mux_module mux_module_inst_2_596(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2105]),.i2(intermediate_reg_1[2104]),.o(intermediate_reg_2[1052]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_597(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2103]),.i2(intermediate_reg_1[2102]),.o(intermediate_reg_2[1051]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_598(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2101]),.i2(intermediate_reg_1[2100]),.o(intermediate_reg_2[1050]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_599(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2099]),.i2(intermediate_reg_1[2098]),.o(intermediate_reg_2[1049])); 
xor_module xor_module_inst_2_600(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2097]),.i2(intermediate_reg_1[2096]),.o(intermediate_reg_2[1048])); 
mux_module mux_module_inst_2_601(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2095]),.i2(intermediate_reg_1[2094]),.o(intermediate_reg_2[1047]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_602(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2093]),.i2(intermediate_reg_1[2092]),.o(intermediate_reg_2[1046]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_603(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2091]),.i2(intermediate_reg_1[2090]),.o(intermediate_reg_2[1045])); 
mux_module mux_module_inst_2_604(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2089]),.i2(intermediate_reg_1[2088]),.o(intermediate_reg_2[1044]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_605(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2087]),.i2(intermediate_reg_1[2086]),.o(intermediate_reg_2[1043]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_606(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2085]),.i2(intermediate_reg_1[2084]),.o(intermediate_reg_2[1042]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_607(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2083]),.i2(intermediate_reg_1[2082]),.o(intermediate_reg_2[1041]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_608(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2081]),.i2(intermediate_reg_1[2080]),.o(intermediate_reg_2[1040])); 
mux_module mux_module_inst_2_609(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2079]),.i2(intermediate_reg_1[2078]),.o(intermediate_reg_2[1039]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_610(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2077]),.i2(intermediate_reg_1[2076]),.o(intermediate_reg_2[1038]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_611(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2075]),.i2(intermediate_reg_1[2074]),.o(intermediate_reg_2[1037])); 
xor_module xor_module_inst_2_612(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2073]),.i2(intermediate_reg_1[2072]),.o(intermediate_reg_2[1036])); 
xor_module xor_module_inst_2_613(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2071]),.i2(intermediate_reg_1[2070]),.o(intermediate_reg_2[1035])); 
mux_module mux_module_inst_2_614(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2069]),.i2(intermediate_reg_1[2068]),.o(intermediate_reg_2[1034]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_615(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2067]),.i2(intermediate_reg_1[2066]),.o(intermediate_reg_2[1033])); 
xor_module xor_module_inst_2_616(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2065]),.i2(intermediate_reg_1[2064]),.o(intermediate_reg_2[1032])); 
mux_module mux_module_inst_2_617(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2063]),.i2(intermediate_reg_1[2062]),.o(intermediate_reg_2[1031]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_618(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2061]),.i2(intermediate_reg_1[2060]),.o(intermediate_reg_2[1030]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_619(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2059]),.i2(intermediate_reg_1[2058]),.o(intermediate_reg_2[1029]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_620(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2057]),.i2(intermediate_reg_1[2056]),.o(intermediate_reg_2[1028])); 
mux_module mux_module_inst_2_621(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2055]),.i2(intermediate_reg_1[2054]),.o(intermediate_reg_2[1027]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_622(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2053]),.i2(intermediate_reg_1[2052]),.o(intermediate_reg_2[1026])); 
mux_module mux_module_inst_2_623(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2051]),.i2(intermediate_reg_1[2050]),.o(intermediate_reg_2[1025]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_624(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2049]),.i2(intermediate_reg_1[2048]),.o(intermediate_reg_2[1024])); 
mux_module mux_module_inst_2_625(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2047]),.i2(intermediate_reg_1[2046]),.o(intermediate_reg_2[1023]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_626(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2045]),.i2(intermediate_reg_1[2044]),.o(intermediate_reg_2[1022])); 
mux_module mux_module_inst_2_627(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2043]),.i2(intermediate_reg_1[2042]),.o(intermediate_reg_2[1021]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_628(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2041]),.i2(intermediate_reg_1[2040]),.o(intermediate_reg_2[1020])); 
mux_module mux_module_inst_2_629(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2039]),.i2(intermediate_reg_1[2038]),.o(intermediate_reg_2[1019]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_630(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2037]),.i2(intermediate_reg_1[2036]),.o(intermediate_reg_2[1018]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_631(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2035]),.i2(intermediate_reg_1[2034]),.o(intermediate_reg_2[1017])); 
mux_module mux_module_inst_2_632(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2033]),.i2(intermediate_reg_1[2032]),.o(intermediate_reg_2[1016]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_633(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2031]),.i2(intermediate_reg_1[2030]),.o(intermediate_reg_2[1015])); 
xor_module xor_module_inst_2_634(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2029]),.i2(intermediate_reg_1[2028]),.o(intermediate_reg_2[1014])); 
xor_module xor_module_inst_2_635(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2027]),.i2(intermediate_reg_1[2026]),.o(intermediate_reg_2[1013])); 
xor_module xor_module_inst_2_636(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2025]),.i2(intermediate_reg_1[2024]),.o(intermediate_reg_2[1012])); 
xor_module xor_module_inst_2_637(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2023]),.i2(intermediate_reg_1[2022]),.o(intermediate_reg_2[1011])); 
xor_module xor_module_inst_2_638(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2021]),.i2(intermediate_reg_1[2020]),.o(intermediate_reg_2[1010])); 
mux_module mux_module_inst_2_639(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2019]),.i2(intermediate_reg_1[2018]),.o(intermediate_reg_2[1009]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_640(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2017]),.i2(intermediate_reg_1[2016]),.o(intermediate_reg_2[1008]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_641(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2015]),.i2(intermediate_reg_1[2014]),.o(intermediate_reg_2[1007])); 
xor_module xor_module_inst_2_642(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2013]),.i2(intermediate_reg_1[2012]),.o(intermediate_reg_2[1006])); 
mux_module mux_module_inst_2_643(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2011]),.i2(intermediate_reg_1[2010]),.o(intermediate_reg_2[1005]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_644(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2009]),.i2(intermediate_reg_1[2008]),.o(intermediate_reg_2[1004]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_645(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2007]),.i2(intermediate_reg_1[2006]),.o(intermediate_reg_2[1003]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_646(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2005]),.i2(intermediate_reg_1[2004]),.o(intermediate_reg_2[1002])); 
mux_module mux_module_inst_2_647(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2003]),.i2(intermediate_reg_1[2002]),.o(intermediate_reg_2[1001]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_648(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2001]),.i2(intermediate_reg_1[2000]),.o(intermediate_reg_2[1000])); 
xor_module xor_module_inst_2_649(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1999]),.i2(intermediate_reg_1[1998]),.o(intermediate_reg_2[999])); 
xor_module xor_module_inst_2_650(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1997]),.i2(intermediate_reg_1[1996]),.o(intermediate_reg_2[998])); 
mux_module mux_module_inst_2_651(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1995]),.i2(intermediate_reg_1[1994]),.o(intermediate_reg_2[997]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_652(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1993]),.i2(intermediate_reg_1[1992]),.o(intermediate_reg_2[996]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_653(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1991]),.i2(intermediate_reg_1[1990]),.o(intermediate_reg_2[995])); 
xor_module xor_module_inst_2_654(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1989]),.i2(intermediate_reg_1[1988]),.o(intermediate_reg_2[994])); 
xor_module xor_module_inst_2_655(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1987]),.i2(intermediate_reg_1[1986]),.o(intermediate_reg_2[993])); 
mux_module mux_module_inst_2_656(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1985]),.i2(intermediate_reg_1[1984]),.o(intermediate_reg_2[992]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_657(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1983]),.i2(intermediate_reg_1[1982]),.o(intermediate_reg_2[991])); 
xor_module xor_module_inst_2_658(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1981]),.i2(intermediate_reg_1[1980]),.o(intermediate_reg_2[990])); 
mux_module mux_module_inst_2_659(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1979]),.i2(intermediate_reg_1[1978]),.o(intermediate_reg_2[989]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_660(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1977]),.i2(intermediate_reg_1[1976]),.o(intermediate_reg_2[988]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_661(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1975]),.i2(intermediate_reg_1[1974]),.o(intermediate_reg_2[987])); 
xor_module xor_module_inst_2_662(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1973]),.i2(intermediate_reg_1[1972]),.o(intermediate_reg_2[986])); 
mux_module mux_module_inst_2_663(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1971]),.i2(intermediate_reg_1[1970]),.o(intermediate_reg_2[985]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_664(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1969]),.i2(intermediate_reg_1[1968]),.o(intermediate_reg_2[984]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_665(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1967]),.i2(intermediate_reg_1[1966]),.o(intermediate_reg_2[983]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_666(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1965]),.i2(intermediate_reg_1[1964]),.o(intermediate_reg_2[982]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_667(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1963]),.i2(intermediate_reg_1[1962]),.o(intermediate_reg_2[981])); 
xor_module xor_module_inst_2_668(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1961]),.i2(intermediate_reg_1[1960]),.o(intermediate_reg_2[980])); 
xor_module xor_module_inst_2_669(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1959]),.i2(intermediate_reg_1[1958]),.o(intermediate_reg_2[979])); 
xor_module xor_module_inst_2_670(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1957]),.i2(intermediate_reg_1[1956]),.o(intermediate_reg_2[978])); 
mux_module mux_module_inst_2_671(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1955]),.i2(intermediate_reg_1[1954]),.o(intermediate_reg_2[977]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_672(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1953]),.i2(intermediate_reg_1[1952]),.o(intermediate_reg_2[976]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_673(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1951]),.i2(intermediate_reg_1[1950]),.o(intermediate_reg_2[975]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_674(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1949]),.i2(intermediate_reg_1[1948]),.o(intermediate_reg_2[974])); 
mux_module mux_module_inst_2_675(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1947]),.i2(intermediate_reg_1[1946]),.o(intermediate_reg_2[973]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_676(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1945]),.i2(intermediate_reg_1[1944]),.o(intermediate_reg_2[972])); 
mux_module mux_module_inst_2_677(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1943]),.i2(intermediate_reg_1[1942]),.o(intermediate_reg_2[971]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_678(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1941]),.i2(intermediate_reg_1[1940]),.o(intermediate_reg_2[970]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_679(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1939]),.i2(intermediate_reg_1[1938]),.o(intermediate_reg_2[969])); 
xor_module xor_module_inst_2_680(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1937]),.i2(intermediate_reg_1[1936]),.o(intermediate_reg_2[968])); 
xor_module xor_module_inst_2_681(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1935]),.i2(intermediate_reg_1[1934]),.o(intermediate_reg_2[967])); 
mux_module mux_module_inst_2_682(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1933]),.i2(intermediate_reg_1[1932]),.o(intermediate_reg_2[966]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_683(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1931]),.i2(intermediate_reg_1[1930]),.o(intermediate_reg_2[965]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_684(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1929]),.i2(intermediate_reg_1[1928]),.o(intermediate_reg_2[964])); 
mux_module mux_module_inst_2_685(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1927]),.i2(intermediate_reg_1[1926]),.o(intermediate_reg_2[963]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_686(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1925]),.i2(intermediate_reg_1[1924]),.o(intermediate_reg_2[962])); 
mux_module mux_module_inst_2_687(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1923]),.i2(intermediate_reg_1[1922]),.o(intermediate_reg_2[961]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_688(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1921]),.i2(intermediate_reg_1[1920]),.o(intermediate_reg_2[960])); 
xor_module xor_module_inst_2_689(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1919]),.i2(intermediate_reg_1[1918]),.o(intermediate_reg_2[959])); 
xor_module xor_module_inst_2_690(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1917]),.i2(intermediate_reg_1[1916]),.o(intermediate_reg_2[958])); 
mux_module mux_module_inst_2_691(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1915]),.i2(intermediate_reg_1[1914]),.o(intermediate_reg_2[957]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_692(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1913]),.i2(intermediate_reg_1[1912]),.o(intermediate_reg_2[956])); 
mux_module mux_module_inst_2_693(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1911]),.i2(intermediate_reg_1[1910]),.o(intermediate_reg_2[955]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_694(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1909]),.i2(intermediate_reg_1[1908]),.o(intermediate_reg_2[954]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_695(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1907]),.i2(intermediate_reg_1[1906]),.o(intermediate_reg_2[953])); 
mux_module mux_module_inst_2_696(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1905]),.i2(intermediate_reg_1[1904]),.o(intermediate_reg_2[952]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_697(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1903]),.i2(intermediate_reg_1[1902]),.o(intermediate_reg_2[951])); 
xor_module xor_module_inst_2_698(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1901]),.i2(intermediate_reg_1[1900]),.o(intermediate_reg_2[950])); 
mux_module mux_module_inst_2_699(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1899]),.i2(intermediate_reg_1[1898]),.o(intermediate_reg_2[949]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_700(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1897]),.i2(intermediate_reg_1[1896]),.o(intermediate_reg_2[948])); 
mux_module mux_module_inst_2_701(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1895]),.i2(intermediate_reg_1[1894]),.o(intermediate_reg_2[947]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_702(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1893]),.i2(intermediate_reg_1[1892]),.o(intermediate_reg_2[946])); 
mux_module mux_module_inst_2_703(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1891]),.i2(intermediate_reg_1[1890]),.o(intermediate_reg_2[945]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_704(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1889]),.i2(intermediate_reg_1[1888]),.o(intermediate_reg_2[944]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_705(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1887]),.i2(intermediate_reg_1[1886]),.o(intermediate_reg_2[943])); 
xor_module xor_module_inst_2_706(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1885]),.i2(intermediate_reg_1[1884]),.o(intermediate_reg_2[942])); 
xor_module xor_module_inst_2_707(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1883]),.i2(intermediate_reg_1[1882]),.o(intermediate_reg_2[941])); 
xor_module xor_module_inst_2_708(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1881]),.i2(intermediate_reg_1[1880]),.o(intermediate_reg_2[940])); 
xor_module xor_module_inst_2_709(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1879]),.i2(intermediate_reg_1[1878]),.o(intermediate_reg_2[939])); 
mux_module mux_module_inst_2_710(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1877]),.i2(intermediate_reg_1[1876]),.o(intermediate_reg_2[938]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_711(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1875]),.i2(intermediate_reg_1[1874]),.o(intermediate_reg_2[937])); 
xor_module xor_module_inst_2_712(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1873]),.i2(intermediate_reg_1[1872]),.o(intermediate_reg_2[936])); 
xor_module xor_module_inst_2_713(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1871]),.i2(intermediate_reg_1[1870]),.o(intermediate_reg_2[935])); 
mux_module mux_module_inst_2_714(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1869]),.i2(intermediate_reg_1[1868]),.o(intermediate_reg_2[934]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_715(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1867]),.i2(intermediate_reg_1[1866]),.o(intermediate_reg_2[933])); 
xor_module xor_module_inst_2_716(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1865]),.i2(intermediate_reg_1[1864]),.o(intermediate_reg_2[932])); 
mux_module mux_module_inst_2_717(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1863]),.i2(intermediate_reg_1[1862]),.o(intermediate_reg_2[931]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_718(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1861]),.i2(intermediate_reg_1[1860]),.o(intermediate_reg_2[930]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_719(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1859]),.i2(intermediate_reg_1[1858]),.o(intermediate_reg_2[929]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_720(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1857]),.i2(intermediate_reg_1[1856]),.o(intermediate_reg_2[928])); 
xor_module xor_module_inst_2_721(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1855]),.i2(intermediate_reg_1[1854]),.o(intermediate_reg_2[927])); 
mux_module mux_module_inst_2_722(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1853]),.i2(intermediate_reg_1[1852]),.o(intermediate_reg_2[926]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_723(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1851]),.i2(intermediate_reg_1[1850]),.o(intermediate_reg_2[925]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_724(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1849]),.i2(intermediate_reg_1[1848]),.o(intermediate_reg_2[924])); 
xor_module xor_module_inst_2_725(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1847]),.i2(intermediate_reg_1[1846]),.o(intermediate_reg_2[923])); 
mux_module mux_module_inst_2_726(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1845]),.i2(intermediate_reg_1[1844]),.o(intermediate_reg_2[922]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_727(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1843]),.i2(intermediate_reg_1[1842]),.o(intermediate_reg_2[921]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_728(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1841]),.i2(intermediate_reg_1[1840]),.o(intermediate_reg_2[920])); 
xor_module xor_module_inst_2_729(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1839]),.i2(intermediate_reg_1[1838]),.o(intermediate_reg_2[919])); 
xor_module xor_module_inst_2_730(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1837]),.i2(intermediate_reg_1[1836]),.o(intermediate_reg_2[918])); 
mux_module mux_module_inst_2_731(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1835]),.i2(intermediate_reg_1[1834]),.o(intermediate_reg_2[917]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_732(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1833]),.i2(intermediate_reg_1[1832]),.o(intermediate_reg_2[916])); 
mux_module mux_module_inst_2_733(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1831]),.i2(intermediate_reg_1[1830]),.o(intermediate_reg_2[915]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_734(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1829]),.i2(intermediate_reg_1[1828]),.o(intermediate_reg_2[914])); 
mux_module mux_module_inst_2_735(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1827]),.i2(intermediate_reg_1[1826]),.o(intermediate_reg_2[913]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_736(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1825]),.i2(intermediate_reg_1[1824]),.o(intermediate_reg_2[912]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_737(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1823]),.i2(intermediate_reg_1[1822]),.o(intermediate_reg_2[911])); 
mux_module mux_module_inst_2_738(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1821]),.i2(intermediate_reg_1[1820]),.o(intermediate_reg_2[910]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_739(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1819]),.i2(intermediate_reg_1[1818]),.o(intermediate_reg_2[909]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_740(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1817]),.i2(intermediate_reg_1[1816]),.o(intermediate_reg_2[908])); 
mux_module mux_module_inst_2_741(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1815]),.i2(intermediate_reg_1[1814]),.o(intermediate_reg_2[907]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_742(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1813]),.i2(intermediate_reg_1[1812]),.o(intermediate_reg_2[906]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_743(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1811]),.i2(intermediate_reg_1[1810]),.o(intermediate_reg_2[905]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_744(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1809]),.i2(intermediate_reg_1[1808]),.o(intermediate_reg_2[904])); 
xor_module xor_module_inst_2_745(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1807]),.i2(intermediate_reg_1[1806]),.o(intermediate_reg_2[903])); 
mux_module mux_module_inst_2_746(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1805]),.i2(intermediate_reg_1[1804]),.o(intermediate_reg_2[902]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_747(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1803]),.i2(intermediate_reg_1[1802]),.o(intermediate_reg_2[901])); 
xor_module xor_module_inst_2_748(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1801]),.i2(intermediate_reg_1[1800]),.o(intermediate_reg_2[900])); 
mux_module mux_module_inst_2_749(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1799]),.i2(intermediate_reg_1[1798]),.o(intermediate_reg_2[899]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_750(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1797]),.i2(intermediate_reg_1[1796]),.o(intermediate_reg_2[898])); 
mux_module mux_module_inst_2_751(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1795]),.i2(intermediate_reg_1[1794]),.o(intermediate_reg_2[897]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_752(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1793]),.i2(intermediate_reg_1[1792]),.o(intermediate_reg_2[896])); 
mux_module mux_module_inst_2_753(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1791]),.i2(intermediate_reg_1[1790]),.o(intermediate_reg_2[895]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_754(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1789]),.i2(intermediate_reg_1[1788]),.o(intermediate_reg_2[894])); 
mux_module mux_module_inst_2_755(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1787]),.i2(intermediate_reg_1[1786]),.o(intermediate_reg_2[893]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_756(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1785]),.i2(intermediate_reg_1[1784]),.o(intermediate_reg_2[892])); 
xor_module xor_module_inst_2_757(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1783]),.i2(intermediate_reg_1[1782]),.o(intermediate_reg_2[891])); 
mux_module mux_module_inst_2_758(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1781]),.i2(intermediate_reg_1[1780]),.o(intermediate_reg_2[890]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_759(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1779]),.i2(intermediate_reg_1[1778]),.o(intermediate_reg_2[889])); 
mux_module mux_module_inst_2_760(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1777]),.i2(intermediate_reg_1[1776]),.o(intermediate_reg_2[888]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_761(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1775]),.i2(intermediate_reg_1[1774]),.o(intermediate_reg_2[887]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_762(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1773]),.i2(intermediate_reg_1[1772]),.o(intermediate_reg_2[886])); 
xor_module xor_module_inst_2_763(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1771]),.i2(intermediate_reg_1[1770]),.o(intermediate_reg_2[885])); 
xor_module xor_module_inst_2_764(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1769]),.i2(intermediate_reg_1[1768]),.o(intermediate_reg_2[884])); 
mux_module mux_module_inst_2_765(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1767]),.i2(intermediate_reg_1[1766]),.o(intermediate_reg_2[883]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_766(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1765]),.i2(intermediate_reg_1[1764]),.o(intermediate_reg_2[882])); 
mux_module mux_module_inst_2_767(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1763]),.i2(intermediate_reg_1[1762]),.o(intermediate_reg_2[881]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_768(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1761]),.i2(intermediate_reg_1[1760]),.o(intermediate_reg_2[880]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_769(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1759]),.i2(intermediate_reg_1[1758]),.o(intermediate_reg_2[879])); 
xor_module xor_module_inst_2_770(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1757]),.i2(intermediate_reg_1[1756]),.o(intermediate_reg_2[878])); 
mux_module mux_module_inst_2_771(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1755]),.i2(intermediate_reg_1[1754]),.o(intermediate_reg_2[877]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_772(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1753]),.i2(intermediate_reg_1[1752]),.o(intermediate_reg_2[876]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_773(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1751]),.i2(intermediate_reg_1[1750]),.o(intermediate_reg_2[875]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_774(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1749]),.i2(intermediate_reg_1[1748]),.o(intermediate_reg_2[874])); 
mux_module mux_module_inst_2_775(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1747]),.i2(intermediate_reg_1[1746]),.o(intermediate_reg_2[873]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_776(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1745]),.i2(intermediate_reg_1[1744]),.o(intermediate_reg_2[872])); 
xor_module xor_module_inst_2_777(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1743]),.i2(intermediate_reg_1[1742]),.o(intermediate_reg_2[871])); 
mux_module mux_module_inst_2_778(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1741]),.i2(intermediate_reg_1[1740]),.o(intermediate_reg_2[870]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_779(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1739]),.i2(intermediate_reg_1[1738]),.o(intermediate_reg_2[869]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_780(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1737]),.i2(intermediate_reg_1[1736]),.o(intermediate_reg_2[868]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_781(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1735]),.i2(intermediate_reg_1[1734]),.o(intermediate_reg_2[867]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_782(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1733]),.i2(intermediate_reg_1[1732]),.o(intermediate_reg_2[866]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_783(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1731]),.i2(intermediate_reg_1[1730]),.o(intermediate_reg_2[865]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_784(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1729]),.i2(intermediate_reg_1[1728]),.o(intermediate_reg_2[864])); 
xor_module xor_module_inst_2_785(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1727]),.i2(intermediate_reg_1[1726]),.o(intermediate_reg_2[863])); 
mux_module mux_module_inst_2_786(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1725]),.i2(intermediate_reg_1[1724]),.o(intermediate_reg_2[862]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_787(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1723]),.i2(intermediate_reg_1[1722]),.o(intermediate_reg_2[861]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_788(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1721]),.i2(intermediate_reg_1[1720]),.o(intermediate_reg_2[860]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_789(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1719]),.i2(intermediate_reg_1[1718]),.o(intermediate_reg_2[859]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_790(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1717]),.i2(intermediate_reg_1[1716]),.o(intermediate_reg_2[858])); 
xor_module xor_module_inst_2_791(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1715]),.i2(intermediate_reg_1[1714]),.o(intermediate_reg_2[857])); 
xor_module xor_module_inst_2_792(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1713]),.i2(intermediate_reg_1[1712]),.o(intermediate_reg_2[856])); 
xor_module xor_module_inst_2_793(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1711]),.i2(intermediate_reg_1[1710]),.o(intermediate_reg_2[855])); 
mux_module mux_module_inst_2_794(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1709]),.i2(intermediate_reg_1[1708]),.o(intermediate_reg_2[854]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_795(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1707]),.i2(intermediate_reg_1[1706]),.o(intermediate_reg_2[853])); 
mux_module mux_module_inst_2_796(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1705]),.i2(intermediate_reg_1[1704]),.o(intermediate_reg_2[852]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_797(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1703]),.i2(intermediate_reg_1[1702]),.o(intermediate_reg_2[851]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_798(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1701]),.i2(intermediate_reg_1[1700]),.o(intermediate_reg_2[850]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_799(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1699]),.i2(intermediate_reg_1[1698]),.o(intermediate_reg_2[849])); 
xor_module xor_module_inst_2_800(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1697]),.i2(intermediate_reg_1[1696]),.o(intermediate_reg_2[848])); 
mux_module mux_module_inst_2_801(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1695]),.i2(intermediate_reg_1[1694]),.o(intermediate_reg_2[847]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_802(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1693]),.i2(intermediate_reg_1[1692]),.o(intermediate_reg_2[846])); 
xor_module xor_module_inst_2_803(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1691]),.i2(intermediate_reg_1[1690]),.o(intermediate_reg_2[845])); 
mux_module mux_module_inst_2_804(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1689]),.i2(intermediate_reg_1[1688]),.o(intermediate_reg_2[844]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_805(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1687]),.i2(intermediate_reg_1[1686]),.o(intermediate_reg_2[843])); 
xor_module xor_module_inst_2_806(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1685]),.i2(intermediate_reg_1[1684]),.o(intermediate_reg_2[842])); 
xor_module xor_module_inst_2_807(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1683]),.i2(intermediate_reg_1[1682]),.o(intermediate_reg_2[841])); 
xor_module xor_module_inst_2_808(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1681]),.i2(intermediate_reg_1[1680]),.o(intermediate_reg_2[840])); 
xor_module xor_module_inst_2_809(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1679]),.i2(intermediate_reg_1[1678]),.o(intermediate_reg_2[839])); 
mux_module mux_module_inst_2_810(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1677]),.i2(intermediate_reg_1[1676]),.o(intermediate_reg_2[838]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_811(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1675]),.i2(intermediate_reg_1[1674]),.o(intermediate_reg_2[837]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_812(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1673]),.i2(intermediate_reg_1[1672]),.o(intermediate_reg_2[836])); 
mux_module mux_module_inst_2_813(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1671]),.i2(intermediate_reg_1[1670]),.o(intermediate_reg_2[835]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_814(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1669]),.i2(intermediate_reg_1[1668]),.o(intermediate_reg_2[834]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_815(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1667]),.i2(intermediate_reg_1[1666]),.o(intermediate_reg_2[833])); 
xor_module xor_module_inst_2_816(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1665]),.i2(intermediate_reg_1[1664]),.o(intermediate_reg_2[832])); 
mux_module mux_module_inst_2_817(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1663]),.i2(intermediate_reg_1[1662]),.o(intermediate_reg_2[831]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_818(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1661]),.i2(intermediate_reg_1[1660]),.o(intermediate_reg_2[830])); 
xor_module xor_module_inst_2_819(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1659]),.i2(intermediate_reg_1[1658]),.o(intermediate_reg_2[829])); 
xor_module xor_module_inst_2_820(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1657]),.i2(intermediate_reg_1[1656]),.o(intermediate_reg_2[828])); 
mux_module mux_module_inst_2_821(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1655]),.i2(intermediate_reg_1[1654]),.o(intermediate_reg_2[827]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_822(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1653]),.i2(intermediate_reg_1[1652]),.o(intermediate_reg_2[826])); 
xor_module xor_module_inst_2_823(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1651]),.i2(intermediate_reg_1[1650]),.o(intermediate_reg_2[825])); 
xor_module xor_module_inst_2_824(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1649]),.i2(intermediate_reg_1[1648]),.o(intermediate_reg_2[824])); 
mux_module mux_module_inst_2_825(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1647]),.i2(intermediate_reg_1[1646]),.o(intermediate_reg_2[823]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_826(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1645]),.i2(intermediate_reg_1[1644]),.o(intermediate_reg_2[822])); 
mux_module mux_module_inst_2_827(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1643]),.i2(intermediate_reg_1[1642]),.o(intermediate_reg_2[821]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_828(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1641]),.i2(intermediate_reg_1[1640]),.o(intermediate_reg_2[820]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_829(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1639]),.i2(intermediate_reg_1[1638]),.o(intermediate_reg_2[819]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_830(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1637]),.i2(intermediate_reg_1[1636]),.o(intermediate_reg_2[818])); 
xor_module xor_module_inst_2_831(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1635]),.i2(intermediate_reg_1[1634]),.o(intermediate_reg_2[817])); 
mux_module mux_module_inst_2_832(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1633]),.i2(intermediate_reg_1[1632]),.o(intermediate_reg_2[816]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_833(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1631]),.i2(intermediate_reg_1[1630]),.o(intermediate_reg_2[815])); 
mux_module mux_module_inst_2_834(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1629]),.i2(intermediate_reg_1[1628]),.o(intermediate_reg_2[814]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_835(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1627]),.i2(intermediate_reg_1[1626]),.o(intermediate_reg_2[813])); 
mux_module mux_module_inst_2_836(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1625]),.i2(intermediate_reg_1[1624]),.o(intermediate_reg_2[812]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_837(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1623]),.i2(intermediate_reg_1[1622]),.o(intermediate_reg_2[811]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_838(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1621]),.i2(intermediate_reg_1[1620]),.o(intermediate_reg_2[810])); 
xor_module xor_module_inst_2_839(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1619]),.i2(intermediate_reg_1[1618]),.o(intermediate_reg_2[809])); 
xor_module xor_module_inst_2_840(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1617]),.i2(intermediate_reg_1[1616]),.o(intermediate_reg_2[808])); 
mux_module mux_module_inst_2_841(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1615]),.i2(intermediate_reg_1[1614]),.o(intermediate_reg_2[807]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_842(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1613]),.i2(intermediate_reg_1[1612]),.o(intermediate_reg_2[806]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_843(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1611]),.i2(intermediate_reg_1[1610]),.o(intermediate_reg_2[805]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_844(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1609]),.i2(intermediate_reg_1[1608]),.o(intermediate_reg_2[804])); 
mux_module mux_module_inst_2_845(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1607]),.i2(intermediate_reg_1[1606]),.o(intermediate_reg_2[803]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_846(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1605]),.i2(intermediate_reg_1[1604]),.o(intermediate_reg_2[802]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_847(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1603]),.i2(intermediate_reg_1[1602]),.o(intermediate_reg_2[801])); 
mux_module mux_module_inst_2_848(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1601]),.i2(intermediate_reg_1[1600]),.o(intermediate_reg_2[800]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_849(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1599]),.i2(intermediate_reg_1[1598]),.o(intermediate_reg_2[799])); 
mux_module mux_module_inst_2_850(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1597]),.i2(intermediate_reg_1[1596]),.o(intermediate_reg_2[798]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_851(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1595]),.i2(intermediate_reg_1[1594]),.o(intermediate_reg_2[797])); 
mux_module mux_module_inst_2_852(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1593]),.i2(intermediate_reg_1[1592]),.o(intermediate_reg_2[796]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_853(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1591]),.i2(intermediate_reg_1[1590]),.o(intermediate_reg_2[795])); 
xor_module xor_module_inst_2_854(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1589]),.i2(intermediate_reg_1[1588]),.o(intermediate_reg_2[794])); 
xor_module xor_module_inst_2_855(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1587]),.i2(intermediate_reg_1[1586]),.o(intermediate_reg_2[793])); 
mux_module mux_module_inst_2_856(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1585]),.i2(intermediate_reg_1[1584]),.o(intermediate_reg_2[792]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_857(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1583]),.i2(intermediate_reg_1[1582]),.o(intermediate_reg_2[791])); 
mux_module mux_module_inst_2_858(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1581]),.i2(intermediate_reg_1[1580]),.o(intermediate_reg_2[790]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_859(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1579]),.i2(intermediate_reg_1[1578]),.o(intermediate_reg_2[789])); 
xor_module xor_module_inst_2_860(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1577]),.i2(intermediate_reg_1[1576]),.o(intermediate_reg_2[788])); 
mux_module mux_module_inst_2_861(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1575]),.i2(intermediate_reg_1[1574]),.o(intermediate_reg_2[787]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_862(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1573]),.i2(intermediate_reg_1[1572]),.o(intermediate_reg_2[786]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_863(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1571]),.i2(intermediate_reg_1[1570]),.o(intermediate_reg_2[785]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_864(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1569]),.i2(intermediate_reg_1[1568]),.o(intermediate_reg_2[784]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_865(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1567]),.i2(intermediate_reg_1[1566]),.o(intermediate_reg_2[783])); 
mux_module mux_module_inst_2_866(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1565]),.i2(intermediate_reg_1[1564]),.o(intermediate_reg_2[782]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_867(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1563]),.i2(intermediate_reg_1[1562]),.o(intermediate_reg_2[781])); 
xor_module xor_module_inst_2_868(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1561]),.i2(intermediate_reg_1[1560]),.o(intermediate_reg_2[780])); 
mux_module mux_module_inst_2_869(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1559]),.i2(intermediate_reg_1[1558]),.o(intermediate_reg_2[779]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_870(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1557]),.i2(intermediate_reg_1[1556]),.o(intermediate_reg_2[778]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_871(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1555]),.i2(intermediate_reg_1[1554]),.o(intermediate_reg_2[777])); 
xor_module xor_module_inst_2_872(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1553]),.i2(intermediate_reg_1[1552]),.o(intermediate_reg_2[776])); 
mux_module mux_module_inst_2_873(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1551]),.i2(intermediate_reg_1[1550]),.o(intermediate_reg_2[775]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_874(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1549]),.i2(intermediate_reg_1[1548]),.o(intermediate_reg_2[774]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_875(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1547]),.i2(intermediate_reg_1[1546]),.o(intermediate_reg_2[773])); 
mux_module mux_module_inst_2_876(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1545]),.i2(intermediate_reg_1[1544]),.o(intermediate_reg_2[772]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_877(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1543]),.i2(intermediate_reg_1[1542]),.o(intermediate_reg_2[771])); 
xor_module xor_module_inst_2_878(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1541]),.i2(intermediate_reg_1[1540]),.o(intermediate_reg_2[770])); 
xor_module xor_module_inst_2_879(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1539]),.i2(intermediate_reg_1[1538]),.o(intermediate_reg_2[769])); 
xor_module xor_module_inst_2_880(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1537]),.i2(intermediate_reg_1[1536]),.o(intermediate_reg_2[768])); 
mux_module mux_module_inst_2_881(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1535]),.i2(intermediate_reg_1[1534]),.o(intermediate_reg_2[767]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_882(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1533]),.i2(intermediate_reg_1[1532]),.o(intermediate_reg_2[766]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_883(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1531]),.i2(intermediate_reg_1[1530]),.o(intermediate_reg_2[765])); 
xor_module xor_module_inst_2_884(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1529]),.i2(intermediate_reg_1[1528]),.o(intermediate_reg_2[764])); 
xor_module xor_module_inst_2_885(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1527]),.i2(intermediate_reg_1[1526]),.o(intermediate_reg_2[763])); 
xor_module xor_module_inst_2_886(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1525]),.i2(intermediate_reg_1[1524]),.o(intermediate_reg_2[762])); 
xor_module xor_module_inst_2_887(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1523]),.i2(intermediate_reg_1[1522]),.o(intermediate_reg_2[761])); 
mux_module mux_module_inst_2_888(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1521]),.i2(intermediate_reg_1[1520]),.o(intermediate_reg_2[760]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_889(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1519]),.i2(intermediate_reg_1[1518]),.o(intermediate_reg_2[759])); 
xor_module xor_module_inst_2_890(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1517]),.i2(intermediate_reg_1[1516]),.o(intermediate_reg_2[758])); 
xor_module xor_module_inst_2_891(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1515]),.i2(intermediate_reg_1[1514]),.o(intermediate_reg_2[757])); 
xor_module xor_module_inst_2_892(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1513]),.i2(intermediate_reg_1[1512]),.o(intermediate_reg_2[756])); 
xor_module xor_module_inst_2_893(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1511]),.i2(intermediate_reg_1[1510]),.o(intermediate_reg_2[755])); 
xor_module xor_module_inst_2_894(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1509]),.i2(intermediate_reg_1[1508]),.o(intermediate_reg_2[754])); 
mux_module mux_module_inst_2_895(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1507]),.i2(intermediate_reg_1[1506]),.o(intermediate_reg_2[753]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_896(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1505]),.i2(intermediate_reg_1[1504]),.o(intermediate_reg_2[752]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_897(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1503]),.i2(intermediate_reg_1[1502]),.o(intermediate_reg_2[751]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_898(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1501]),.i2(intermediate_reg_1[1500]),.o(intermediate_reg_2[750]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_899(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1499]),.i2(intermediate_reg_1[1498]),.o(intermediate_reg_2[749]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_900(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1497]),.i2(intermediate_reg_1[1496]),.o(intermediate_reg_2[748]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_901(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1495]),.i2(intermediate_reg_1[1494]),.o(intermediate_reg_2[747])); 
mux_module mux_module_inst_2_902(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1493]),.i2(intermediate_reg_1[1492]),.o(intermediate_reg_2[746]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_903(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1491]),.i2(intermediate_reg_1[1490]),.o(intermediate_reg_2[745]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_904(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1489]),.i2(intermediate_reg_1[1488]),.o(intermediate_reg_2[744])); 
xor_module xor_module_inst_2_905(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1487]),.i2(intermediate_reg_1[1486]),.o(intermediate_reg_2[743])); 
mux_module mux_module_inst_2_906(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1485]),.i2(intermediate_reg_1[1484]),.o(intermediate_reg_2[742]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_907(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1483]),.i2(intermediate_reg_1[1482]),.o(intermediate_reg_2[741])); 
xor_module xor_module_inst_2_908(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1481]),.i2(intermediate_reg_1[1480]),.o(intermediate_reg_2[740])); 
mux_module mux_module_inst_2_909(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1479]),.i2(intermediate_reg_1[1478]),.o(intermediate_reg_2[739]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_910(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1477]),.i2(intermediate_reg_1[1476]),.o(intermediate_reg_2[738]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_911(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1475]),.i2(intermediate_reg_1[1474]),.o(intermediate_reg_2[737]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_912(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1473]),.i2(intermediate_reg_1[1472]),.o(intermediate_reg_2[736])); 
xor_module xor_module_inst_2_913(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1471]),.i2(intermediate_reg_1[1470]),.o(intermediate_reg_2[735])); 
mux_module mux_module_inst_2_914(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1469]),.i2(intermediate_reg_1[1468]),.o(intermediate_reg_2[734]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_915(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1467]),.i2(intermediate_reg_1[1466]),.o(intermediate_reg_2[733]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_916(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1465]),.i2(intermediate_reg_1[1464]),.o(intermediate_reg_2[732]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_917(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1463]),.i2(intermediate_reg_1[1462]),.o(intermediate_reg_2[731])); 
xor_module xor_module_inst_2_918(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1461]),.i2(intermediate_reg_1[1460]),.o(intermediate_reg_2[730])); 
mux_module mux_module_inst_2_919(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1459]),.i2(intermediate_reg_1[1458]),.o(intermediate_reg_2[729]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_920(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1457]),.i2(intermediate_reg_1[1456]),.o(intermediate_reg_2[728])); 
xor_module xor_module_inst_2_921(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1455]),.i2(intermediate_reg_1[1454]),.o(intermediate_reg_2[727])); 
mux_module mux_module_inst_2_922(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1453]),.i2(intermediate_reg_1[1452]),.o(intermediate_reg_2[726]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_923(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1451]),.i2(intermediate_reg_1[1450]),.o(intermediate_reg_2[725]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_924(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1449]),.i2(intermediate_reg_1[1448]),.o(intermediate_reg_2[724])); 
mux_module mux_module_inst_2_925(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1447]),.i2(intermediate_reg_1[1446]),.o(intermediate_reg_2[723]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_926(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1445]),.i2(intermediate_reg_1[1444]),.o(intermediate_reg_2[722]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_927(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1443]),.i2(intermediate_reg_1[1442]),.o(intermediate_reg_2[721])); 
xor_module xor_module_inst_2_928(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1441]),.i2(intermediate_reg_1[1440]),.o(intermediate_reg_2[720])); 
mux_module mux_module_inst_2_929(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1439]),.i2(intermediate_reg_1[1438]),.o(intermediate_reg_2[719]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_930(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1437]),.i2(intermediate_reg_1[1436]),.o(intermediate_reg_2[718]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_931(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1435]),.i2(intermediate_reg_1[1434]),.o(intermediate_reg_2[717])); 
mux_module mux_module_inst_2_932(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1433]),.i2(intermediate_reg_1[1432]),.o(intermediate_reg_2[716]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_933(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1431]),.i2(intermediate_reg_1[1430]),.o(intermediate_reg_2[715]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_934(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1429]),.i2(intermediate_reg_1[1428]),.o(intermediate_reg_2[714])); 
mux_module mux_module_inst_2_935(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1427]),.i2(intermediate_reg_1[1426]),.o(intermediate_reg_2[713]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_936(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1425]),.i2(intermediate_reg_1[1424]),.o(intermediate_reg_2[712])); 
mux_module mux_module_inst_2_937(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1423]),.i2(intermediate_reg_1[1422]),.o(intermediate_reg_2[711]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_938(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1421]),.i2(intermediate_reg_1[1420]),.o(intermediate_reg_2[710]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_939(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1419]),.i2(intermediate_reg_1[1418]),.o(intermediate_reg_2[709])); 
mux_module mux_module_inst_2_940(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1417]),.i2(intermediate_reg_1[1416]),.o(intermediate_reg_2[708]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_941(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1415]),.i2(intermediate_reg_1[1414]),.o(intermediate_reg_2[707]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_942(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1413]),.i2(intermediate_reg_1[1412]),.o(intermediate_reg_2[706]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_943(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1411]),.i2(intermediate_reg_1[1410]),.o(intermediate_reg_2[705]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_944(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1409]),.i2(intermediate_reg_1[1408]),.o(intermediate_reg_2[704]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_945(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1407]),.i2(intermediate_reg_1[1406]),.o(intermediate_reg_2[703])); 
xor_module xor_module_inst_2_946(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1405]),.i2(intermediate_reg_1[1404]),.o(intermediate_reg_2[702])); 
xor_module xor_module_inst_2_947(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1403]),.i2(intermediate_reg_1[1402]),.o(intermediate_reg_2[701])); 
xor_module xor_module_inst_2_948(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1401]),.i2(intermediate_reg_1[1400]),.o(intermediate_reg_2[700])); 
xor_module xor_module_inst_2_949(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1399]),.i2(intermediate_reg_1[1398]),.o(intermediate_reg_2[699])); 
xor_module xor_module_inst_2_950(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1397]),.i2(intermediate_reg_1[1396]),.o(intermediate_reg_2[698])); 
mux_module mux_module_inst_2_951(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1395]),.i2(intermediate_reg_1[1394]),.o(intermediate_reg_2[697]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_952(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1393]),.i2(intermediate_reg_1[1392]),.o(intermediate_reg_2[696]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_953(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1391]),.i2(intermediate_reg_1[1390]),.o(intermediate_reg_2[695]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_954(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1389]),.i2(intermediate_reg_1[1388]),.o(intermediate_reg_2[694])); 
xor_module xor_module_inst_2_955(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1387]),.i2(intermediate_reg_1[1386]),.o(intermediate_reg_2[693])); 
xor_module xor_module_inst_2_956(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1385]),.i2(intermediate_reg_1[1384]),.o(intermediate_reg_2[692])); 
xor_module xor_module_inst_2_957(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1383]),.i2(intermediate_reg_1[1382]),.o(intermediate_reg_2[691])); 
xor_module xor_module_inst_2_958(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1381]),.i2(intermediate_reg_1[1380]),.o(intermediate_reg_2[690])); 
mux_module mux_module_inst_2_959(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1379]),.i2(intermediate_reg_1[1378]),.o(intermediate_reg_2[689]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_960(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1377]),.i2(intermediate_reg_1[1376]),.o(intermediate_reg_2[688]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_961(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1375]),.i2(intermediate_reg_1[1374]),.o(intermediate_reg_2[687])); 
xor_module xor_module_inst_2_962(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1373]),.i2(intermediate_reg_1[1372]),.o(intermediate_reg_2[686])); 
mux_module mux_module_inst_2_963(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1371]),.i2(intermediate_reg_1[1370]),.o(intermediate_reg_2[685]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_964(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1369]),.i2(intermediate_reg_1[1368]),.o(intermediate_reg_2[684]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_965(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1367]),.i2(intermediate_reg_1[1366]),.o(intermediate_reg_2[683]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_966(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1365]),.i2(intermediate_reg_1[1364]),.o(intermediate_reg_2[682]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_967(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1363]),.i2(intermediate_reg_1[1362]),.o(intermediate_reg_2[681]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_968(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1361]),.i2(intermediate_reg_1[1360]),.o(intermediate_reg_2[680])); 
xor_module xor_module_inst_2_969(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1359]),.i2(intermediate_reg_1[1358]),.o(intermediate_reg_2[679])); 
xor_module xor_module_inst_2_970(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1357]),.i2(intermediate_reg_1[1356]),.o(intermediate_reg_2[678])); 
mux_module mux_module_inst_2_971(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1355]),.i2(intermediate_reg_1[1354]),.o(intermediate_reg_2[677]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_972(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1353]),.i2(intermediate_reg_1[1352]),.o(intermediate_reg_2[676]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_973(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1351]),.i2(intermediate_reg_1[1350]),.o(intermediate_reg_2[675])); 
xor_module xor_module_inst_2_974(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1349]),.i2(intermediate_reg_1[1348]),.o(intermediate_reg_2[674])); 
mux_module mux_module_inst_2_975(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1347]),.i2(intermediate_reg_1[1346]),.o(intermediate_reg_2[673]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_976(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1345]),.i2(intermediate_reg_1[1344]),.o(intermediate_reg_2[672]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_977(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1343]),.i2(intermediate_reg_1[1342]),.o(intermediate_reg_2[671]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_978(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1341]),.i2(intermediate_reg_1[1340]),.o(intermediate_reg_2[670])); 
xor_module xor_module_inst_2_979(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1339]),.i2(intermediate_reg_1[1338]),.o(intermediate_reg_2[669])); 
mux_module mux_module_inst_2_980(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1337]),.i2(intermediate_reg_1[1336]),.o(intermediate_reg_2[668]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_981(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1335]),.i2(intermediate_reg_1[1334]),.o(intermediate_reg_2[667]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_982(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1333]),.i2(intermediate_reg_1[1332]),.o(intermediate_reg_2[666])); 
mux_module mux_module_inst_2_983(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1331]),.i2(intermediate_reg_1[1330]),.o(intermediate_reg_2[665]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_984(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1329]),.i2(intermediate_reg_1[1328]),.o(intermediate_reg_2[664])); 
xor_module xor_module_inst_2_985(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1327]),.i2(intermediate_reg_1[1326]),.o(intermediate_reg_2[663])); 
mux_module mux_module_inst_2_986(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1325]),.i2(intermediate_reg_1[1324]),.o(intermediate_reg_2[662]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_987(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1323]),.i2(intermediate_reg_1[1322]),.o(intermediate_reg_2[661]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_988(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1321]),.i2(intermediate_reg_1[1320]),.o(intermediate_reg_2[660]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_989(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1319]),.i2(intermediate_reg_1[1318]),.o(intermediate_reg_2[659]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_990(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1317]),.i2(intermediate_reg_1[1316]),.o(intermediate_reg_2[658])); 
xor_module xor_module_inst_2_991(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1315]),.i2(intermediate_reg_1[1314]),.o(intermediate_reg_2[657])); 
mux_module mux_module_inst_2_992(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1313]),.i2(intermediate_reg_1[1312]),.o(intermediate_reg_2[656]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_993(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1311]),.i2(intermediate_reg_1[1310]),.o(intermediate_reg_2[655])); 
mux_module mux_module_inst_2_994(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1309]),.i2(intermediate_reg_1[1308]),.o(intermediate_reg_2[654]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_995(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1307]),.i2(intermediate_reg_1[1306]),.o(intermediate_reg_2[653]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_996(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1305]),.i2(intermediate_reg_1[1304]),.o(intermediate_reg_2[652])); 
xor_module xor_module_inst_2_997(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1303]),.i2(intermediate_reg_1[1302]),.o(intermediate_reg_2[651])); 
mux_module mux_module_inst_2_998(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1301]),.i2(intermediate_reg_1[1300]),.o(intermediate_reg_2[650]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_999(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1299]),.i2(intermediate_reg_1[1298]),.o(intermediate_reg_2[649])); 
mux_module mux_module_inst_2_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1297]),.i2(intermediate_reg_1[1296]),.o(intermediate_reg_2[648]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1295]),.i2(intermediate_reg_1[1294]),.o(intermediate_reg_2[647]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1293]),.i2(intermediate_reg_1[1292]),.o(intermediate_reg_2[646]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1291]),.i2(intermediate_reg_1[1290]),.o(intermediate_reg_2[645]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1289]),.i2(intermediate_reg_1[1288]),.o(intermediate_reg_2[644])); 
mux_module mux_module_inst_2_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1287]),.i2(intermediate_reg_1[1286]),.o(intermediate_reg_2[643]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1285]),.i2(intermediate_reg_1[1284]),.o(intermediate_reg_2[642]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1283]),.i2(intermediate_reg_1[1282]),.o(intermediate_reg_2[641])); 
mux_module mux_module_inst_2_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1281]),.i2(intermediate_reg_1[1280]),.o(intermediate_reg_2[640]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1279]),.i2(intermediate_reg_1[1278]),.o(intermediate_reg_2[639]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1277]),.i2(intermediate_reg_1[1276]),.o(intermediate_reg_2[638])); 
mux_module mux_module_inst_2_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1275]),.i2(intermediate_reg_1[1274]),.o(intermediate_reg_2[637]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1273]),.i2(intermediate_reg_1[1272]),.o(intermediate_reg_2[636])); 
xor_module xor_module_inst_2_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1271]),.i2(intermediate_reg_1[1270]),.o(intermediate_reg_2[635])); 
xor_module xor_module_inst_2_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1269]),.i2(intermediate_reg_1[1268]),.o(intermediate_reg_2[634])); 
xor_module xor_module_inst_2_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1267]),.i2(intermediate_reg_1[1266]),.o(intermediate_reg_2[633])); 
mux_module mux_module_inst_2_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1265]),.i2(intermediate_reg_1[1264]),.o(intermediate_reg_2[632]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1263]),.i2(intermediate_reg_1[1262]),.o(intermediate_reg_2[631])); 
xor_module xor_module_inst_2_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1261]),.i2(intermediate_reg_1[1260]),.o(intermediate_reg_2[630])); 
mux_module mux_module_inst_2_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1259]),.i2(intermediate_reg_1[1258]),.o(intermediate_reg_2[629]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1257]),.i2(intermediate_reg_1[1256]),.o(intermediate_reg_2[628])); 
xor_module xor_module_inst_2_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1255]),.i2(intermediate_reg_1[1254]),.o(intermediate_reg_2[627])); 
mux_module mux_module_inst_2_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1253]),.i2(intermediate_reg_1[1252]),.o(intermediate_reg_2[626]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1251]),.i2(intermediate_reg_1[1250]),.o(intermediate_reg_2[625]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1249]),.i2(intermediate_reg_1[1248]),.o(intermediate_reg_2[624]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1247]),.i2(intermediate_reg_1[1246]),.o(intermediate_reg_2[623]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1245]),.i2(intermediate_reg_1[1244]),.o(intermediate_reg_2[622])); 
xor_module xor_module_inst_2_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1243]),.i2(intermediate_reg_1[1242]),.o(intermediate_reg_2[621])); 
xor_module xor_module_inst_2_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1241]),.i2(intermediate_reg_1[1240]),.o(intermediate_reg_2[620])); 
mux_module mux_module_inst_2_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1239]),.i2(intermediate_reg_1[1238]),.o(intermediate_reg_2[619]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1237]),.i2(intermediate_reg_1[1236]),.o(intermediate_reg_2[618]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1235]),.i2(intermediate_reg_1[1234]),.o(intermediate_reg_2[617]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1233]),.i2(intermediate_reg_1[1232]),.o(intermediate_reg_2[616]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1231]),.i2(intermediate_reg_1[1230]),.o(intermediate_reg_2[615])); 
mux_module mux_module_inst_2_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1229]),.i2(intermediate_reg_1[1228]),.o(intermediate_reg_2[614]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1227]),.i2(intermediate_reg_1[1226]),.o(intermediate_reg_2[613])); 
xor_module xor_module_inst_2_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1225]),.i2(intermediate_reg_1[1224]),.o(intermediate_reg_2[612])); 
mux_module mux_module_inst_2_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1223]),.i2(intermediate_reg_1[1222]),.o(intermediate_reg_2[611]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1221]),.i2(intermediate_reg_1[1220]),.o(intermediate_reg_2[610]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1219]),.i2(intermediate_reg_1[1218]),.o(intermediate_reg_2[609])); 
mux_module mux_module_inst_2_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1217]),.i2(intermediate_reg_1[1216]),.o(intermediate_reg_2[608]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1215]),.i2(intermediate_reg_1[1214]),.o(intermediate_reg_2[607])); 
mux_module mux_module_inst_2_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1213]),.i2(intermediate_reg_1[1212]),.o(intermediate_reg_2[606]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1211]),.i2(intermediate_reg_1[1210]),.o(intermediate_reg_2[605]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1209]),.i2(intermediate_reg_1[1208]),.o(intermediate_reg_2[604]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1207]),.i2(intermediate_reg_1[1206]),.o(intermediate_reg_2[603]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1205]),.i2(intermediate_reg_1[1204]),.o(intermediate_reg_2[602])); 
mux_module mux_module_inst_2_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1203]),.i2(intermediate_reg_1[1202]),.o(intermediate_reg_2[601]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1201]),.i2(intermediate_reg_1[1200]),.o(intermediate_reg_2[600])); 
xor_module xor_module_inst_2_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1199]),.i2(intermediate_reg_1[1198]),.o(intermediate_reg_2[599])); 
mux_module mux_module_inst_2_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1197]),.i2(intermediate_reg_1[1196]),.o(intermediate_reg_2[598]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1195]),.i2(intermediate_reg_1[1194]),.o(intermediate_reg_2[597]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1193]),.i2(intermediate_reg_1[1192]),.o(intermediate_reg_2[596]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1191]),.i2(intermediate_reg_1[1190]),.o(intermediate_reg_2[595]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1189]),.i2(intermediate_reg_1[1188]),.o(intermediate_reg_2[594])); 
xor_module xor_module_inst_2_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1187]),.i2(intermediate_reg_1[1186]),.o(intermediate_reg_2[593])); 
xor_module xor_module_inst_2_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1185]),.i2(intermediate_reg_1[1184]),.o(intermediate_reg_2[592])); 
mux_module mux_module_inst_2_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1183]),.i2(intermediate_reg_1[1182]),.o(intermediate_reg_2[591]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1181]),.i2(intermediate_reg_1[1180]),.o(intermediate_reg_2[590]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1179]),.i2(intermediate_reg_1[1178]),.o(intermediate_reg_2[589])); 
xor_module xor_module_inst_2_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1177]),.i2(intermediate_reg_1[1176]),.o(intermediate_reg_2[588])); 
xor_module xor_module_inst_2_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1175]),.i2(intermediate_reg_1[1174]),.o(intermediate_reg_2[587])); 
mux_module mux_module_inst_2_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1173]),.i2(intermediate_reg_1[1172]),.o(intermediate_reg_2[586]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1171]),.i2(intermediate_reg_1[1170]),.o(intermediate_reg_2[585]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1169]),.i2(intermediate_reg_1[1168]),.o(intermediate_reg_2[584]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1167]),.i2(intermediate_reg_1[1166]),.o(intermediate_reg_2[583])); 
xor_module xor_module_inst_2_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1165]),.i2(intermediate_reg_1[1164]),.o(intermediate_reg_2[582])); 
mux_module mux_module_inst_2_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1163]),.i2(intermediate_reg_1[1162]),.o(intermediate_reg_2[581]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1161]),.i2(intermediate_reg_1[1160]),.o(intermediate_reg_2[580]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1159]),.i2(intermediate_reg_1[1158]),.o(intermediate_reg_2[579]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1157]),.i2(intermediate_reg_1[1156]),.o(intermediate_reg_2[578])); 
mux_module mux_module_inst_2_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1155]),.i2(intermediate_reg_1[1154]),.o(intermediate_reg_2[577]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1153]),.i2(intermediate_reg_1[1152]),.o(intermediate_reg_2[576]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1151]),.i2(intermediate_reg_1[1150]),.o(intermediate_reg_2[575])); 
xor_module xor_module_inst_2_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1149]),.i2(intermediate_reg_1[1148]),.o(intermediate_reg_2[574])); 
xor_module xor_module_inst_2_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1147]),.i2(intermediate_reg_1[1146]),.o(intermediate_reg_2[573])); 
mux_module mux_module_inst_2_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1145]),.i2(intermediate_reg_1[1144]),.o(intermediate_reg_2[572]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1143]),.i2(intermediate_reg_1[1142]),.o(intermediate_reg_2[571]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1141]),.i2(intermediate_reg_1[1140]),.o(intermediate_reg_2[570]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1139]),.i2(intermediate_reg_1[1138]),.o(intermediate_reg_2[569])); 
mux_module mux_module_inst_2_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1137]),.i2(intermediate_reg_1[1136]),.o(intermediate_reg_2[568]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1135]),.i2(intermediate_reg_1[1134]),.o(intermediate_reg_2[567]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1133]),.i2(intermediate_reg_1[1132]),.o(intermediate_reg_2[566])); 
xor_module xor_module_inst_2_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1131]),.i2(intermediate_reg_1[1130]),.o(intermediate_reg_2[565])); 
xor_module xor_module_inst_2_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1129]),.i2(intermediate_reg_1[1128]),.o(intermediate_reg_2[564])); 
mux_module mux_module_inst_2_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1127]),.i2(intermediate_reg_1[1126]),.o(intermediate_reg_2[563]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1125]),.i2(intermediate_reg_1[1124]),.o(intermediate_reg_2[562]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1123]),.i2(intermediate_reg_1[1122]),.o(intermediate_reg_2[561]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1121]),.i2(intermediate_reg_1[1120]),.o(intermediate_reg_2[560]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1119]),.i2(intermediate_reg_1[1118]),.o(intermediate_reg_2[559]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1117]),.i2(intermediate_reg_1[1116]),.o(intermediate_reg_2[558])); 
mux_module mux_module_inst_2_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1115]),.i2(intermediate_reg_1[1114]),.o(intermediate_reg_2[557]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1113]),.i2(intermediate_reg_1[1112]),.o(intermediate_reg_2[556]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1111]),.i2(intermediate_reg_1[1110]),.o(intermediate_reg_2[555]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1109]),.i2(intermediate_reg_1[1108]),.o(intermediate_reg_2[554])); 
xor_module xor_module_inst_2_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1107]),.i2(intermediate_reg_1[1106]),.o(intermediate_reg_2[553])); 
mux_module mux_module_inst_2_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1105]),.i2(intermediate_reg_1[1104]),.o(intermediate_reg_2[552]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1103]),.i2(intermediate_reg_1[1102]),.o(intermediate_reg_2[551])); 
mux_module mux_module_inst_2_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1101]),.i2(intermediate_reg_1[1100]),.o(intermediate_reg_2[550]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1099]),.i2(intermediate_reg_1[1098]),.o(intermediate_reg_2[549]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1097]),.i2(intermediate_reg_1[1096]),.o(intermediate_reg_2[548])); 
mux_module mux_module_inst_2_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1095]),.i2(intermediate_reg_1[1094]),.o(intermediate_reg_2[547]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1093]),.i2(intermediate_reg_1[1092]),.o(intermediate_reg_2[546]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1091]),.i2(intermediate_reg_1[1090]),.o(intermediate_reg_2[545]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1089]),.i2(intermediate_reg_1[1088]),.o(intermediate_reg_2[544]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1087]),.i2(intermediate_reg_1[1086]),.o(intermediate_reg_2[543]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1085]),.i2(intermediate_reg_1[1084]),.o(intermediate_reg_2[542])); 
mux_module mux_module_inst_2_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1083]),.i2(intermediate_reg_1[1082]),.o(intermediate_reg_2[541]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1081]),.i2(intermediate_reg_1[1080]),.o(intermediate_reg_2[540])); 
xor_module xor_module_inst_2_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1079]),.i2(intermediate_reg_1[1078]),.o(intermediate_reg_2[539])); 
xor_module xor_module_inst_2_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1077]),.i2(intermediate_reg_1[1076]),.o(intermediate_reg_2[538])); 
xor_module xor_module_inst_2_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1075]),.i2(intermediate_reg_1[1074]),.o(intermediate_reg_2[537])); 
xor_module xor_module_inst_2_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1073]),.i2(intermediate_reg_1[1072]),.o(intermediate_reg_2[536])); 
xor_module xor_module_inst_2_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1071]),.i2(intermediate_reg_1[1070]),.o(intermediate_reg_2[535])); 
mux_module mux_module_inst_2_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1069]),.i2(intermediate_reg_1[1068]),.o(intermediate_reg_2[534]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1067]),.i2(intermediate_reg_1[1066]),.o(intermediate_reg_2[533])); 
xor_module xor_module_inst_2_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1065]),.i2(intermediate_reg_1[1064]),.o(intermediate_reg_2[532])); 
mux_module mux_module_inst_2_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1063]),.i2(intermediate_reg_1[1062]),.o(intermediate_reg_2[531]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1061]),.i2(intermediate_reg_1[1060]),.o(intermediate_reg_2[530])); 
xor_module xor_module_inst_2_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1059]),.i2(intermediate_reg_1[1058]),.o(intermediate_reg_2[529])); 
mux_module mux_module_inst_2_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1057]),.i2(intermediate_reg_1[1056]),.o(intermediate_reg_2[528]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1055]),.i2(intermediate_reg_1[1054]),.o(intermediate_reg_2[527])); 
xor_module xor_module_inst_2_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1053]),.i2(intermediate_reg_1[1052]),.o(intermediate_reg_2[526])); 
mux_module mux_module_inst_2_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1051]),.i2(intermediate_reg_1[1050]),.o(intermediate_reg_2[525]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1049]),.i2(intermediate_reg_1[1048]),.o(intermediate_reg_2[524]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1047]),.i2(intermediate_reg_1[1046]),.o(intermediate_reg_2[523]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1045]),.i2(intermediate_reg_1[1044]),.o(intermediate_reg_2[522])); 
mux_module mux_module_inst_2_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1043]),.i2(intermediate_reg_1[1042]),.o(intermediate_reg_2[521]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1041]),.i2(intermediate_reg_1[1040]),.o(intermediate_reg_2[520]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1039]),.i2(intermediate_reg_1[1038]),.o(intermediate_reg_2[519]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1037]),.i2(intermediate_reg_1[1036]),.o(intermediate_reg_2[518])); 
xor_module xor_module_inst_2_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1035]),.i2(intermediate_reg_1[1034]),.o(intermediate_reg_2[517])); 
xor_module xor_module_inst_2_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1033]),.i2(intermediate_reg_1[1032]),.o(intermediate_reg_2[516])); 
mux_module mux_module_inst_2_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1031]),.i2(intermediate_reg_1[1030]),.o(intermediate_reg_2[515]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1029]),.i2(intermediate_reg_1[1028]),.o(intermediate_reg_2[514])); 
xor_module xor_module_inst_2_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1027]),.i2(intermediate_reg_1[1026]),.o(intermediate_reg_2[513])); 
mux_module mux_module_inst_2_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1025]),.i2(intermediate_reg_1[1024]),.o(intermediate_reg_2[512]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1023]),.i2(intermediate_reg_1[1022]),.o(intermediate_reg_2[511]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1021]),.i2(intermediate_reg_1[1020]),.o(intermediate_reg_2[510])); 
xor_module xor_module_inst_2_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1019]),.i2(intermediate_reg_1[1018]),.o(intermediate_reg_2[509])); 
xor_module xor_module_inst_2_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1017]),.i2(intermediate_reg_1[1016]),.o(intermediate_reg_2[508])); 
mux_module mux_module_inst_2_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1015]),.i2(intermediate_reg_1[1014]),.o(intermediate_reg_2[507]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1013]),.i2(intermediate_reg_1[1012]),.o(intermediate_reg_2[506])); 
mux_module mux_module_inst_2_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1011]),.i2(intermediate_reg_1[1010]),.o(intermediate_reg_2[505]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1009]),.i2(intermediate_reg_1[1008]),.o(intermediate_reg_2[504]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1007]),.i2(intermediate_reg_1[1006]),.o(intermediate_reg_2[503])); 
mux_module mux_module_inst_2_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1005]),.i2(intermediate_reg_1[1004]),.o(intermediate_reg_2[502]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1003]),.i2(intermediate_reg_1[1002]),.o(intermediate_reg_2[501])); 
mux_module mux_module_inst_2_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1001]),.i2(intermediate_reg_1[1000]),.o(intermediate_reg_2[500]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[999]),.i2(intermediate_reg_1[998]),.o(intermediate_reg_2[499])); 
mux_module mux_module_inst_2_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[997]),.i2(intermediate_reg_1[996]),.o(intermediate_reg_2[498]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[995]),.i2(intermediate_reg_1[994]),.o(intermediate_reg_2[497]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[993]),.i2(intermediate_reg_1[992]),.o(intermediate_reg_2[496]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[991]),.i2(intermediate_reg_1[990]),.o(intermediate_reg_2[495]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[989]),.i2(intermediate_reg_1[988]),.o(intermediate_reg_2[494])); 
xor_module xor_module_inst_2_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[987]),.i2(intermediate_reg_1[986]),.o(intermediate_reg_2[493])); 
xor_module xor_module_inst_2_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[985]),.i2(intermediate_reg_1[984]),.o(intermediate_reg_2[492])); 
xor_module xor_module_inst_2_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[983]),.i2(intermediate_reg_1[982]),.o(intermediate_reg_2[491])); 
xor_module xor_module_inst_2_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[981]),.i2(intermediate_reg_1[980]),.o(intermediate_reg_2[490])); 
mux_module mux_module_inst_2_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[979]),.i2(intermediate_reg_1[978]),.o(intermediate_reg_2[489]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[977]),.i2(intermediate_reg_1[976]),.o(intermediate_reg_2[488]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[975]),.i2(intermediate_reg_1[974]),.o(intermediate_reg_2[487]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[973]),.i2(intermediate_reg_1[972]),.o(intermediate_reg_2[486]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[971]),.i2(intermediate_reg_1[970]),.o(intermediate_reg_2[485])); 
mux_module mux_module_inst_2_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[969]),.i2(intermediate_reg_1[968]),.o(intermediate_reg_2[484]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[967]),.i2(intermediate_reg_1[966]),.o(intermediate_reg_2[483]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[965]),.i2(intermediate_reg_1[964]),.o(intermediate_reg_2[482])); 
xor_module xor_module_inst_2_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[963]),.i2(intermediate_reg_1[962]),.o(intermediate_reg_2[481])); 
xor_module xor_module_inst_2_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[961]),.i2(intermediate_reg_1[960]),.o(intermediate_reg_2[480])); 
xor_module xor_module_inst_2_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479])); 
xor_module xor_module_inst_2_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478])); 
mux_module mux_module_inst_2_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472])); 
mux_module mux_module_inst_2_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466])); 
xor_module xor_module_inst_2_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465])); 
xor_module xor_module_inst_2_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464])); 
mux_module mux_module_inst_2_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454])); 
xor_module xor_module_inst_2_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453])); 
xor_module xor_module_inst_2_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452])); 
mux_module mux_module_inst_2_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448])); 
xor_module xor_module_inst_2_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447])); 
mux_module mux_module_inst_2_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445])); 
xor_module xor_module_inst_2_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444])); 
mux_module mux_module_inst_2_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438])); 
mux_module mux_module_inst_2_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436])); 
mux_module mux_module_inst_2_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434])); 
xor_module xor_module_inst_2_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433])); 
xor_module xor_module_inst_2_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432])); 
mux_module mux_module_inst_2_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430])); 
mux_module mux_module_inst_2_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428])); 
mux_module mux_module_inst_2_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426])); 
xor_module xor_module_inst_2_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425])); 
xor_module xor_module_inst_2_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424])); 
mux_module mux_module_inst_2_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422])); 
xor_module xor_module_inst_2_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421])); 
mux_module mux_module_inst_2_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418])); 
xor_module xor_module_inst_2_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417])); 
mux_module mux_module_inst_2_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415])); 
xor_module xor_module_inst_2_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414])); 
mux_module mux_module_inst_2_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410])); 
xor_module xor_module_inst_2_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409])); 
xor_module xor_module_inst_2_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408])); 
xor_module xor_module_inst_2_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407])); 
xor_module xor_module_inst_2_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406])); 
mux_module mux_module_inst_2_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401])); 
mux_module mux_module_inst_2_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398])); 
xor_module xor_module_inst_2_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397])); 
mux_module mux_module_inst_2_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395])); 
xor_module xor_module_inst_2_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394])); 
xor_module xor_module_inst_2_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393])); 
xor_module xor_module_inst_2_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392])); 
mux_module mux_module_inst_2_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390])); 
mux_module mux_module_inst_2_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387])); 
mux_module mux_module_inst_2_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384])); 
mux_module mux_module_inst_2_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381])); 
xor_module xor_module_inst_2_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380])); 
xor_module xor_module_inst_2_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379])); 
mux_module mux_module_inst_2_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375])); 
xor_module xor_module_inst_2_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374])); 
mux_module mux_module_inst_2_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372])); 
mux_module mux_module_inst_2_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370])); 
xor_module xor_module_inst_2_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369])); 
mux_module mux_module_inst_2_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366])); 
mux_module mux_module_inst_2_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364])); 
xor_module xor_module_inst_2_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363])); 
mux_module mux_module_inst_2_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361])); 
xor_module xor_module_inst_2_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360])); 
xor_module xor_module_inst_2_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359])); 
xor_module xor_module_inst_2_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358])); 
xor_module xor_module_inst_2_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357])); 
mux_module mux_module_inst_2_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355])); 
mux_module mux_module_inst_2_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349])); 
xor_module xor_module_inst_2_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348])); 
xor_module xor_module_inst_2_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347])); 
mux_module mux_module_inst_2_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343])); 
mux_module mux_module_inst_2_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340])); 
xor_module xor_module_inst_2_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339])); 
xor_module xor_module_inst_2_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338])); 
xor_module xor_module_inst_2_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337])); 
xor_module xor_module_inst_2_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336])); 
xor_module xor_module_inst_2_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335])); 
mux_module mux_module_inst_2_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332])); 
xor_module xor_module_inst_2_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331])); 
mux_module mux_module_inst_2_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329])); 
xor_module xor_module_inst_2_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328])); 
xor_module xor_module_inst_2_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327])); 
xor_module xor_module_inst_2_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326])); 
xor_module xor_module_inst_2_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325])); 
mux_module mux_module_inst_2_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323])); 
mux_module mux_module_inst_2_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320])); 
xor_module xor_module_inst_2_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319])); 
mux_module mux_module_inst_2_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316])); 
xor_module xor_module_inst_2_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315])); 
mux_module mux_module_inst_2_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311])); 
mux_module mux_module_inst_2_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308])); 
xor_module xor_module_inst_2_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307])); 
xor_module xor_module_inst_2_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306])); 
mux_module mux_module_inst_2_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304])); 
mux_module mux_module_inst_2_1345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300])); 
xor_module xor_module_inst_2_1349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299])); 
xor_module xor_module_inst_2_1350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298])); 
mux_module mux_module_inst_2_1351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293])); 
xor_module xor_module_inst_2_1356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292])); 
xor_module xor_module_inst_2_1357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291])); 
xor_module xor_module_inst_2_1358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290])); 
mux_module mux_module_inst_2_1359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286])); 
xor_module xor_module_inst_2_1363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
xor_module xor_module_inst_2_1364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284])); 
xor_module xor_module_inst_2_1365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
xor_module xor_module_inst_2_1366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282])); 
mux_module mux_module_inst_2_1367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279])); 
xor_module xor_module_inst_2_1370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278])); 
mux_module mux_module_inst_2_1371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272])); 
mux_module mux_module_inst_2_1377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270])); 
xor_module xor_module_inst_2_1379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269])); 
mux_module mux_module_inst_2_1380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266])); 
xor_module xor_module_inst_2_1383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265])); 
mux_module mux_module_inst_2_1384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263])); 
mux_module mux_module_inst_2_1386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261])); 
xor_module xor_module_inst_2_1388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260])); 
mux_module mux_module_inst_2_1389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258])); 
mux_module mux_module_inst_2_1391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
mux_module mux_module_inst_2_1393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254])); 
xor_module xor_module_inst_2_1395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253])); 
xor_module xor_module_inst_2_1396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252])); 
xor_module xor_module_inst_2_1397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251])); 
xor_module xor_module_inst_2_1398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250])); 
mux_module mux_module_inst_2_1399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
xor_module xor_module_inst_2_1404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244])); 
xor_module xor_module_inst_2_1405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243])); 
xor_module xor_module_inst_2_1406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242])); 
mux_module mux_module_inst_2_1407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235])); 
xor_module xor_module_inst_2_1414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
xor_module xor_module_inst_2_1415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233])); 
xor_module xor_module_inst_2_1416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232])); 
xor_module xor_module_inst_2_1417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231])); 
mux_module mux_module_inst_2_1418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226])); 
mux_module mux_module_inst_2_1423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224])); 
xor_module xor_module_inst_2_1425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223])); 
xor_module xor_module_inst_2_1426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
xor_module xor_module_inst_2_1427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221])); 
xor_module xor_module_inst_2_1428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220])); 
xor_module xor_module_inst_2_1429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219])); 
mux_module mux_module_inst_2_1430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217])); 
xor_module xor_module_inst_2_1432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216])); 
mux_module mux_module_inst_2_1433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214])); 
xor_module xor_module_inst_2_1435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
mux_module mux_module_inst_2_1436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211])); 
xor_module xor_module_inst_2_1438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
mux_module mux_module_inst_2_1439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208])); 
mux_module mux_module_inst_2_1441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
mux_module mux_module_inst_2_1443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197])); 
mux_module mux_module_inst_2_1452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193])); 
xor_module xor_module_inst_2_1456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
xor_module xor_module_inst_2_1457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
mux_module mux_module_inst_2_1458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187])); 
mux_module mux_module_inst_2_1462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
xor_module xor_module_inst_2_1465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183])); 
mux_module mux_module_inst_2_1466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177])); 
mux_module mux_module_inst_2_1472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
xor_module xor_module_inst_2_1476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
mux_module mux_module_inst_2_1477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
mux_module mux_module_inst_2_1479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168])); 
mux_module mux_module_inst_2_1481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162])); 
xor_module xor_module_inst_2_1487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161])); 
mux_module mux_module_inst_2_1488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
mux_module mux_module_inst_2_1490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156])); 
xor_module xor_module_inst_2_1493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155])); 
mux_module mux_module_inst_2_1494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152])); 
xor_module xor_module_inst_2_1497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151])); 
xor_module xor_module_inst_2_1498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
xor_module xor_module_inst_2_1499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
mux_module mux_module_inst_2_1500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147])); 
mux_module mux_module_inst_2_1502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145])); 
xor_module xor_module_inst_2_1504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144])); 
mux_module mux_module_inst_2_1505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142])); 
xor_module xor_module_inst_2_1507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141])); 
mux_module mux_module_inst_2_1508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137])); 
xor_module xor_module_inst_2_1512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136])); 
mux_module mux_module_inst_2_1513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1514(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
mux_module mux_module_inst_2_1515(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1516(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1517(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1518(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1519(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129])); 
xor_module xor_module_inst_2_1520(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
xor_module xor_module_inst_2_1521(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127])); 
mux_module mux_module_inst_2_1522(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1523(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
xor_module xor_module_inst_2_1524(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124])); 
xor_module xor_module_inst_2_1525(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123])); 
xor_module xor_module_inst_2_1526(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122])); 
xor_module xor_module_inst_2_1527(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121])); 
mux_module mux_module_inst_2_1528(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1529(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1530(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1531(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117])); 
mux_module mux_module_inst_2_1532(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1533(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115])); 
xor_module xor_module_inst_2_1534(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114])); 
mux_module mux_module_inst_2_1535(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1536(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
mux_module mux_module_inst_2_1537(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1538(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
mux_module mux_module_inst_2_1539(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1540(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108])); 
mux_module mux_module_inst_2_1541(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1542(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
xor_module xor_module_inst_2_1543(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105])); 
mux_module mux_module_inst_2_1544(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1545(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103])); 
xor_module xor_module_inst_2_1546(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102])); 
xor_module xor_module_inst_2_1547(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101])); 
xor_module xor_module_inst_2_1548(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100])); 
mux_module mux_module_inst_2_1549(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1550(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1551(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1552(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96])); 
xor_module xor_module_inst_2_1553(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95])); 
mux_module mux_module_inst_2_1554(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1555(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
xor_module xor_module_inst_2_1556(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92])); 
mux_module mux_module_inst_2_1557(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1558(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90])); 
xor_module xor_module_inst_2_1559(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89])); 
xor_module xor_module_inst_2_1560(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88])); 
xor_module xor_module_inst_2_1561(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
xor_module xor_module_inst_2_1562(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86])); 
xor_module xor_module_inst_2_1563(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
mux_module mux_module_inst_2_1564(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1565(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83])); 
xor_module xor_module_inst_2_1566(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82])); 
mux_module mux_module_inst_2_1567(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1568(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80])); 
xor_module xor_module_inst_2_1569(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79])); 
xor_module xor_module_inst_2_1570(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78])); 
xor_module xor_module_inst_2_1571(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77])); 
xor_module xor_module_inst_2_1572(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76])); 
mux_module mux_module_inst_2_1573(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1574(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74])); 
xor_module xor_module_inst_2_1575(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73])); 
mux_module mux_module_inst_2_1576(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1577(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71])); 
xor_module xor_module_inst_2_1578(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
mux_module mux_module_inst_2_1579(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1580(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68])); 
mux_module mux_module_inst_2_1581(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1582(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1583(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1584(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1585(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63])); 
xor_module xor_module_inst_2_1586(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
xor_module xor_module_inst_2_1587(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
xor_module xor_module_inst_2_1588(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60])); 
mux_module mux_module_inst_2_1589(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1590(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58])); 
xor_module xor_module_inst_2_1591(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57])); 
mux_module mux_module_inst_2_1592(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1593(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1594(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1595(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
xor_module xor_module_inst_2_1596(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
xor_module xor_module_inst_2_1597(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51])); 
mux_module mux_module_inst_2_1598(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1599(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
xor_module xor_module_inst_2_1600(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48])); 
xor_module xor_module_inst_2_1601(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47])); 
xor_module xor_module_inst_2_1602(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46])); 
mux_module mux_module_inst_2_1603(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1604(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1605(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43])); 
xor_module xor_module_inst_2_1606(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42])); 
xor_module xor_module_inst_2_1607(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41])); 
xor_module xor_module_inst_2_1608(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40])); 
mux_module mux_module_inst_2_1609(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1610(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38])); 
mux_module mux_module_inst_2_1611(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1612(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36])); 
xor_module xor_module_inst_2_1613(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35])); 
xor_module xor_module_inst_2_1614(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34])); 
mux_module mux_module_inst_2_1615(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1616(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32])); 
xor_module xor_module_inst_2_1617(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31])); 
xor_module xor_module_inst_2_1618(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30])); 
mux_module mux_module_inst_2_1619(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1620(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1621(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27])); 
mux_module mux_module_inst_2_1622(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1623(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1624(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24])); 
xor_module xor_module_inst_2_1625(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23])); 
xor_module xor_module_inst_2_1626(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22])); 
mux_module mux_module_inst_2_1627(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1628(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20])); 
mux_module mux_module_inst_2_1629(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1630(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1631(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17])); 
xor_module xor_module_inst_2_1632(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16])); 
xor_module xor_module_inst_2_1633(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15])); 
mux_module mux_module_inst_2_1634(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1635(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1636(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1637(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1638(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1639(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9])); 
xor_module xor_module_inst_2_1640(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8])); 
mux_module mux_module_inst_2_1641(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1642(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6])); 
mux_module mux_module_inst_2_1643(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1644(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
xor_module xor_module_inst_2_1645(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
mux_module mux_module_inst_2_1646(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1647(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1648(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0]),.sel(intermediate_reg_1[0])); 
wire [1647:0]intermediate_wire_3; 
assign intermediate_wire_3[1647] = intermediate_reg_2[1648]^intermediate_reg_2[1647] ; 
assign intermediate_wire_3[1646:0] = intermediate_reg_2[1646:0] ; 
wire [823:0]intermediate_reg_3; 
 
xor_module xor_module_inst_3_0(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1647]),.i2(intermediate_wire_3[1646]),.o(intermediate_reg_3[823])); 
xor_module xor_module_inst_3_1(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1645]),.i2(intermediate_wire_3[1644]),.o(intermediate_reg_3[822])); 
mux_module mux_module_inst_3_2(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1643]),.i2(intermediate_wire_3[1642]),.o(intermediate_reg_3[821]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_3(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1641]),.i2(intermediate_wire_3[1640]),.o(intermediate_reg_3[820])); 
mux_module mux_module_inst_3_4(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1639]),.i2(intermediate_wire_3[1638]),.o(intermediate_reg_3[819]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_5(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1637]),.i2(intermediate_wire_3[1636]),.o(intermediate_reg_3[818])); 
mux_module mux_module_inst_3_6(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1635]),.i2(intermediate_wire_3[1634]),.o(intermediate_reg_3[817]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_7(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1633]),.i2(intermediate_wire_3[1632]),.o(intermediate_reg_3[816]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_8(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1631]),.i2(intermediate_wire_3[1630]),.o(intermediate_reg_3[815])); 
mux_module mux_module_inst_3_9(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1629]),.i2(intermediate_wire_3[1628]),.o(intermediate_reg_3[814]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_10(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1627]),.i2(intermediate_wire_3[1626]),.o(intermediate_reg_3[813])); 
mux_module mux_module_inst_3_11(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1625]),.i2(intermediate_wire_3[1624]),.o(intermediate_reg_3[812]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_12(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1623]),.i2(intermediate_wire_3[1622]),.o(intermediate_reg_3[811])); 
xor_module xor_module_inst_3_13(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1621]),.i2(intermediate_wire_3[1620]),.o(intermediate_reg_3[810])); 
mux_module mux_module_inst_3_14(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1619]),.i2(intermediate_wire_3[1618]),.o(intermediate_reg_3[809]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_15(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1617]),.i2(intermediate_wire_3[1616]),.o(intermediate_reg_3[808]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_16(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1615]),.i2(intermediate_wire_3[1614]),.o(intermediate_reg_3[807])); 
mux_module mux_module_inst_3_17(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1613]),.i2(intermediate_wire_3[1612]),.o(intermediate_reg_3[806]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_18(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1611]),.i2(intermediate_wire_3[1610]),.o(intermediate_reg_3[805])); 
xor_module xor_module_inst_3_19(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1609]),.i2(intermediate_wire_3[1608]),.o(intermediate_reg_3[804])); 
xor_module xor_module_inst_3_20(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1607]),.i2(intermediate_wire_3[1606]),.o(intermediate_reg_3[803])); 
xor_module xor_module_inst_3_21(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1605]),.i2(intermediate_wire_3[1604]),.o(intermediate_reg_3[802])); 
mux_module mux_module_inst_3_22(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1603]),.i2(intermediate_wire_3[1602]),.o(intermediate_reg_3[801]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_23(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1601]),.i2(intermediate_wire_3[1600]),.o(intermediate_reg_3[800])); 
xor_module xor_module_inst_3_24(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1599]),.i2(intermediate_wire_3[1598]),.o(intermediate_reg_3[799])); 
xor_module xor_module_inst_3_25(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1597]),.i2(intermediate_wire_3[1596]),.o(intermediate_reg_3[798])); 
xor_module xor_module_inst_3_26(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1595]),.i2(intermediate_wire_3[1594]),.o(intermediate_reg_3[797])); 
mux_module mux_module_inst_3_27(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1593]),.i2(intermediate_wire_3[1592]),.o(intermediate_reg_3[796]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_28(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1591]),.i2(intermediate_wire_3[1590]),.o(intermediate_reg_3[795])); 
xor_module xor_module_inst_3_29(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1589]),.i2(intermediate_wire_3[1588]),.o(intermediate_reg_3[794])); 
mux_module mux_module_inst_3_30(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1587]),.i2(intermediate_wire_3[1586]),.o(intermediate_reg_3[793]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_31(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1585]),.i2(intermediate_wire_3[1584]),.o(intermediate_reg_3[792])); 
xor_module xor_module_inst_3_32(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1583]),.i2(intermediate_wire_3[1582]),.o(intermediate_reg_3[791])); 
xor_module xor_module_inst_3_33(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1581]),.i2(intermediate_wire_3[1580]),.o(intermediate_reg_3[790])); 
mux_module mux_module_inst_3_34(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1579]),.i2(intermediate_wire_3[1578]),.o(intermediate_reg_3[789]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_35(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1577]),.i2(intermediate_wire_3[1576]),.o(intermediate_reg_3[788]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_36(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1575]),.i2(intermediate_wire_3[1574]),.o(intermediate_reg_3[787])); 
xor_module xor_module_inst_3_37(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1573]),.i2(intermediate_wire_3[1572]),.o(intermediate_reg_3[786])); 
xor_module xor_module_inst_3_38(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1571]),.i2(intermediate_wire_3[1570]),.o(intermediate_reg_3[785])); 
xor_module xor_module_inst_3_39(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1569]),.i2(intermediate_wire_3[1568]),.o(intermediate_reg_3[784])); 
mux_module mux_module_inst_3_40(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1567]),.i2(intermediate_wire_3[1566]),.o(intermediate_reg_3[783]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_41(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1565]),.i2(intermediate_wire_3[1564]),.o(intermediate_reg_3[782])); 
xor_module xor_module_inst_3_42(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1563]),.i2(intermediate_wire_3[1562]),.o(intermediate_reg_3[781])); 
xor_module xor_module_inst_3_43(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1561]),.i2(intermediate_wire_3[1560]),.o(intermediate_reg_3[780])); 
mux_module mux_module_inst_3_44(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1559]),.i2(intermediate_wire_3[1558]),.o(intermediate_reg_3[779]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_45(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1557]),.i2(intermediate_wire_3[1556]),.o(intermediate_reg_3[778])); 
mux_module mux_module_inst_3_46(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1555]),.i2(intermediate_wire_3[1554]),.o(intermediate_reg_3[777]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_47(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1553]),.i2(intermediate_wire_3[1552]),.o(intermediate_reg_3[776]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_48(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1551]),.i2(intermediate_wire_3[1550]),.o(intermediate_reg_3[775])); 
mux_module mux_module_inst_3_49(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1549]),.i2(intermediate_wire_3[1548]),.o(intermediate_reg_3[774]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_50(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1547]),.i2(intermediate_wire_3[1546]),.o(intermediate_reg_3[773])); 
mux_module mux_module_inst_3_51(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1545]),.i2(intermediate_wire_3[1544]),.o(intermediate_reg_3[772]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_52(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1543]),.i2(intermediate_wire_3[1542]),.o(intermediate_reg_3[771])); 
xor_module xor_module_inst_3_53(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1541]),.i2(intermediate_wire_3[1540]),.o(intermediate_reg_3[770])); 
mux_module mux_module_inst_3_54(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1539]),.i2(intermediate_wire_3[1538]),.o(intermediate_reg_3[769]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_55(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1537]),.i2(intermediate_wire_3[1536]),.o(intermediate_reg_3[768]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_56(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1535]),.i2(intermediate_wire_3[1534]),.o(intermediate_reg_3[767])); 
mux_module mux_module_inst_3_57(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1533]),.i2(intermediate_wire_3[1532]),.o(intermediate_reg_3[766]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_58(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1531]),.i2(intermediate_wire_3[1530]),.o(intermediate_reg_3[765]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_59(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1529]),.i2(intermediate_wire_3[1528]),.o(intermediate_reg_3[764]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_60(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1527]),.i2(intermediate_wire_3[1526]),.o(intermediate_reg_3[763]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_61(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1525]),.i2(intermediate_wire_3[1524]),.o(intermediate_reg_3[762]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_62(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1523]),.i2(intermediate_wire_3[1522]),.o(intermediate_reg_3[761])); 
mux_module mux_module_inst_3_63(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1521]),.i2(intermediate_wire_3[1520]),.o(intermediate_reg_3[760]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_64(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1519]),.i2(intermediate_wire_3[1518]),.o(intermediate_reg_3[759]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_65(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1517]),.i2(intermediate_wire_3[1516]),.o(intermediate_reg_3[758])); 
mux_module mux_module_inst_3_66(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1515]),.i2(intermediate_wire_3[1514]),.o(intermediate_reg_3[757]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_67(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1513]),.i2(intermediate_wire_3[1512]),.o(intermediate_reg_3[756]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_68(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1511]),.i2(intermediate_wire_3[1510]),.o(intermediate_reg_3[755])); 
xor_module xor_module_inst_3_69(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1509]),.i2(intermediate_wire_3[1508]),.o(intermediate_reg_3[754])); 
xor_module xor_module_inst_3_70(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1507]),.i2(intermediate_wire_3[1506]),.o(intermediate_reg_3[753])); 
mux_module mux_module_inst_3_71(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1505]),.i2(intermediate_wire_3[1504]),.o(intermediate_reg_3[752]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_72(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1503]),.i2(intermediate_wire_3[1502]),.o(intermediate_reg_3[751]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_73(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1501]),.i2(intermediate_wire_3[1500]),.o(intermediate_reg_3[750]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_74(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1499]),.i2(intermediate_wire_3[1498]),.o(intermediate_reg_3[749]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_75(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1497]),.i2(intermediate_wire_3[1496]),.o(intermediate_reg_3[748])); 
xor_module xor_module_inst_3_76(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1495]),.i2(intermediate_wire_3[1494]),.o(intermediate_reg_3[747])); 
xor_module xor_module_inst_3_77(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1493]),.i2(intermediate_wire_3[1492]),.o(intermediate_reg_3[746])); 
mux_module mux_module_inst_3_78(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1491]),.i2(intermediate_wire_3[1490]),.o(intermediate_reg_3[745]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_79(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1489]),.i2(intermediate_wire_3[1488]),.o(intermediate_reg_3[744])); 
xor_module xor_module_inst_3_80(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1487]),.i2(intermediate_wire_3[1486]),.o(intermediate_reg_3[743])); 
mux_module mux_module_inst_3_81(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1485]),.i2(intermediate_wire_3[1484]),.o(intermediate_reg_3[742]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_82(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1483]),.i2(intermediate_wire_3[1482]),.o(intermediate_reg_3[741])); 
xor_module xor_module_inst_3_83(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1481]),.i2(intermediate_wire_3[1480]),.o(intermediate_reg_3[740])); 
mux_module mux_module_inst_3_84(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1479]),.i2(intermediate_wire_3[1478]),.o(intermediate_reg_3[739]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_85(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1477]),.i2(intermediate_wire_3[1476]),.o(intermediate_reg_3[738]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_86(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1475]),.i2(intermediate_wire_3[1474]),.o(intermediate_reg_3[737]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_87(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1473]),.i2(intermediate_wire_3[1472]),.o(intermediate_reg_3[736])); 
mux_module mux_module_inst_3_88(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1471]),.i2(intermediate_wire_3[1470]),.o(intermediate_reg_3[735]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_89(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1469]),.i2(intermediate_wire_3[1468]),.o(intermediate_reg_3[734]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_90(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1467]),.i2(intermediate_wire_3[1466]),.o(intermediate_reg_3[733]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_91(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1465]),.i2(intermediate_wire_3[1464]),.o(intermediate_reg_3[732])); 
xor_module xor_module_inst_3_92(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1463]),.i2(intermediate_wire_3[1462]),.o(intermediate_reg_3[731])); 
mux_module mux_module_inst_3_93(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1461]),.i2(intermediate_wire_3[1460]),.o(intermediate_reg_3[730]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_94(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1459]),.i2(intermediate_wire_3[1458]),.o(intermediate_reg_3[729])); 
xor_module xor_module_inst_3_95(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1457]),.i2(intermediate_wire_3[1456]),.o(intermediate_reg_3[728])); 
xor_module xor_module_inst_3_96(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1455]),.i2(intermediate_wire_3[1454]),.o(intermediate_reg_3[727])); 
xor_module xor_module_inst_3_97(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1453]),.i2(intermediate_wire_3[1452]),.o(intermediate_reg_3[726])); 
mux_module mux_module_inst_3_98(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1451]),.i2(intermediate_wire_3[1450]),.o(intermediate_reg_3[725]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_99(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1449]),.i2(intermediate_wire_3[1448]),.o(intermediate_reg_3[724])); 
mux_module mux_module_inst_3_100(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1447]),.i2(intermediate_wire_3[1446]),.o(intermediate_reg_3[723]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_101(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1445]),.i2(intermediate_wire_3[1444]),.o(intermediate_reg_3[722]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_102(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1443]),.i2(intermediate_wire_3[1442]),.o(intermediate_reg_3[721])); 
mux_module mux_module_inst_3_103(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1441]),.i2(intermediate_wire_3[1440]),.o(intermediate_reg_3[720]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_104(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1439]),.i2(intermediate_wire_3[1438]),.o(intermediate_reg_3[719])); 
mux_module mux_module_inst_3_105(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1437]),.i2(intermediate_wire_3[1436]),.o(intermediate_reg_3[718]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_106(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1435]),.i2(intermediate_wire_3[1434]),.o(intermediate_reg_3[717])); 
xor_module xor_module_inst_3_107(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1433]),.i2(intermediate_wire_3[1432]),.o(intermediate_reg_3[716])); 
mux_module mux_module_inst_3_108(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1431]),.i2(intermediate_wire_3[1430]),.o(intermediate_reg_3[715]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_109(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1429]),.i2(intermediate_wire_3[1428]),.o(intermediate_reg_3[714])); 
mux_module mux_module_inst_3_110(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1427]),.i2(intermediate_wire_3[1426]),.o(intermediate_reg_3[713]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_111(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1425]),.i2(intermediate_wire_3[1424]),.o(intermediate_reg_3[712]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_112(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1423]),.i2(intermediate_wire_3[1422]),.o(intermediate_reg_3[711]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_113(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1421]),.i2(intermediate_wire_3[1420]),.o(intermediate_reg_3[710]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_114(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1419]),.i2(intermediate_wire_3[1418]),.o(intermediate_reg_3[709])); 
xor_module xor_module_inst_3_115(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1417]),.i2(intermediate_wire_3[1416]),.o(intermediate_reg_3[708])); 
xor_module xor_module_inst_3_116(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1415]),.i2(intermediate_wire_3[1414]),.o(intermediate_reg_3[707])); 
mux_module mux_module_inst_3_117(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1413]),.i2(intermediate_wire_3[1412]),.o(intermediate_reg_3[706]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_118(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1411]),.i2(intermediate_wire_3[1410]),.o(intermediate_reg_3[705]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_119(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1409]),.i2(intermediate_wire_3[1408]),.o(intermediate_reg_3[704])); 
mux_module mux_module_inst_3_120(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1407]),.i2(intermediate_wire_3[1406]),.o(intermediate_reg_3[703]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_121(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1405]),.i2(intermediate_wire_3[1404]),.o(intermediate_reg_3[702])); 
xor_module xor_module_inst_3_122(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1403]),.i2(intermediate_wire_3[1402]),.o(intermediate_reg_3[701])); 
xor_module xor_module_inst_3_123(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1401]),.i2(intermediate_wire_3[1400]),.o(intermediate_reg_3[700])); 
mux_module mux_module_inst_3_124(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1399]),.i2(intermediate_wire_3[1398]),.o(intermediate_reg_3[699]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_125(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1397]),.i2(intermediate_wire_3[1396]),.o(intermediate_reg_3[698])); 
mux_module mux_module_inst_3_126(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1395]),.i2(intermediate_wire_3[1394]),.o(intermediate_reg_3[697]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_127(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1393]),.i2(intermediate_wire_3[1392]),.o(intermediate_reg_3[696]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_128(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1391]),.i2(intermediate_wire_3[1390]),.o(intermediate_reg_3[695])); 
xor_module xor_module_inst_3_129(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1389]),.i2(intermediate_wire_3[1388]),.o(intermediate_reg_3[694])); 
mux_module mux_module_inst_3_130(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1387]),.i2(intermediate_wire_3[1386]),.o(intermediate_reg_3[693]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_131(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1385]),.i2(intermediate_wire_3[1384]),.o(intermediate_reg_3[692]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_132(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1383]),.i2(intermediate_wire_3[1382]),.o(intermediate_reg_3[691])); 
mux_module mux_module_inst_3_133(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1381]),.i2(intermediate_wire_3[1380]),.o(intermediate_reg_3[690]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_134(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1379]),.i2(intermediate_wire_3[1378]),.o(intermediate_reg_3[689])); 
mux_module mux_module_inst_3_135(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1377]),.i2(intermediate_wire_3[1376]),.o(intermediate_reg_3[688]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_136(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1375]),.i2(intermediate_wire_3[1374]),.o(intermediate_reg_3[687])); 
xor_module xor_module_inst_3_137(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1373]),.i2(intermediate_wire_3[1372]),.o(intermediate_reg_3[686])); 
mux_module mux_module_inst_3_138(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1371]),.i2(intermediate_wire_3[1370]),.o(intermediate_reg_3[685]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_139(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1369]),.i2(intermediate_wire_3[1368]),.o(intermediate_reg_3[684])); 
xor_module xor_module_inst_3_140(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1367]),.i2(intermediate_wire_3[1366]),.o(intermediate_reg_3[683])); 
xor_module xor_module_inst_3_141(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1365]),.i2(intermediate_wire_3[1364]),.o(intermediate_reg_3[682])); 
mux_module mux_module_inst_3_142(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1363]),.i2(intermediate_wire_3[1362]),.o(intermediate_reg_3[681]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_143(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1361]),.i2(intermediate_wire_3[1360]),.o(intermediate_reg_3[680]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_144(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1359]),.i2(intermediate_wire_3[1358]),.o(intermediate_reg_3[679])); 
xor_module xor_module_inst_3_145(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1357]),.i2(intermediate_wire_3[1356]),.o(intermediate_reg_3[678])); 
mux_module mux_module_inst_3_146(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1355]),.i2(intermediate_wire_3[1354]),.o(intermediate_reg_3[677]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_147(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1353]),.i2(intermediate_wire_3[1352]),.o(intermediate_reg_3[676]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_148(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1351]),.i2(intermediate_wire_3[1350]),.o(intermediate_reg_3[675]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_149(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1349]),.i2(intermediate_wire_3[1348]),.o(intermediate_reg_3[674]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_150(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1347]),.i2(intermediate_wire_3[1346]),.o(intermediate_reg_3[673]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_151(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1345]),.i2(intermediate_wire_3[1344]),.o(intermediate_reg_3[672]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_152(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1343]),.i2(intermediate_wire_3[1342]),.o(intermediate_reg_3[671])); 
mux_module mux_module_inst_3_153(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1341]),.i2(intermediate_wire_3[1340]),.o(intermediate_reg_3[670]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_154(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1339]),.i2(intermediate_wire_3[1338]),.o(intermediate_reg_3[669])); 
xor_module xor_module_inst_3_155(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1337]),.i2(intermediate_wire_3[1336]),.o(intermediate_reg_3[668])); 
mux_module mux_module_inst_3_156(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1335]),.i2(intermediate_wire_3[1334]),.o(intermediate_reg_3[667]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_157(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1333]),.i2(intermediate_wire_3[1332]),.o(intermediate_reg_3[666])); 
mux_module mux_module_inst_3_158(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1331]),.i2(intermediate_wire_3[1330]),.o(intermediate_reg_3[665]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_159(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1329]),.i2(intermediate_wire_3[1328]),.o(intermediate_reg_3[664]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_160(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1327]),.i2(intermediate_wire_3[1326]),.o(intermediate_reg_3[663])); 
xor_module xor_module_inst_3_161(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1325]),.i2(intermediate_wire_3[1324]),.o(intermediate_reg_3[662])); 
mux_module mux_module_inst_3_162(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1323]),.i2(intermediate_wire_3[1322]),.o(intermediate_reg_3[661]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_163(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1321]),.i2(intermediate_wire_3[1320]),.o(intermediate_reg_3[660]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_164(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1319]),.i2(intermediate_wire_3[1318]),.o(intermediate_reg_3[659])); 
mux_module mux_module_inst_3_165(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1317]),.i2(intermediate_wire_3[1316]),.o(intermediate_reg_3[658]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_166(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1315]),.i2(intermediate_wire_3[1314]),.o(intermediate_reg_3[657]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_167(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1313]),.i2(intermediate_wire_3[1312]),.o(intermediate_reg_3[656]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_168(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1311]),.i2(intermediate_wire_3[1310]),.o(intermediate_reg_3[655])); 
xor_module xor_module_inst_3_169(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1309]),.i2(intermediate_wire_3[1308]),.o(intermediate_reg_3[654])); 
xor_module xor_module_inst_3_170(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1307]),.i2(intermediate_wire_3[1306]),.o(intermediate_reg_3[653])); 
mux_module mux_module_inst_3_171(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1305]),.i2(intermediate_wire_3[1304]),.o(intermediate_reg_3[652]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_172(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1303]),.i2(intermediate_wire_3[1302]),.o(intermediate_reg_3[651]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_173(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1301]),.i2(intermediate_wire_3[1300]),.o(intermediate_reg_3[650]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_174(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1299]),.i2(intermediate_wire_3[1298]),.o(intermediate_reg_3[649])); 
mux_module mux_module_inst_3_175(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1297]),.i2(intermediate_wire_3[1296]),.o(intermediate_reg_3[648]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_176(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1295]),.i2(intermediate_wire_3[1294]),.o(intermediate_reg_3[647])); 
xor_module xor_module_inst_3_177(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1293]),.i2(intermediate_wire_3[1292]),.o(intermediate_reg_3[646])); 
xor_module xor_module_inst_3_178(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1291]),.i2(intermediate_wire_3[1290]),.o(intermediate_reg_3[645])); 
mux_module mux_module_inst_3_179(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1289]),.i2(intermediate_wire_3[1288]),.o(intermediate_reg_3[644]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_180(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1287]),.i2(intermediate_wire_3[1286]),.o(intermediate_reg_3[643])); 
mux_module mux_module_inst_3_181(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1285]),.i2(intermediate_wire_3[1284]),.o(intermediate_reg_3[642]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_182(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1283]),.i2(intermediate_wire_3[1282]),.o(intermediate_reg_3[641]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_183(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1281]),.i2(intermediate_wire_3[1280]),.o(intermediate_reg_3[640]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_184(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1279]),.i2(intermediate_wire_3[1278]),.o(intermediate_reg_3[639]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_185(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1277]),.i2(intermediate_wire_3[1276]),.o(intermediate_reg_3[638]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_186(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1275]),.i2(intermediate_wire_3[1274]),.o(intermediate_reg_3[637])); 
xor_module xor_module_inst_3_187(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1273]),.i2(intermediate_wire_3[1272]),.o(intermediate_reg_3[636])); 
mux_module mux_module_inst_3_188(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1271]),.i2(intermediate_wire_3[1270]),.o(intermediate_reg_3[635]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_189(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1269]),.i2(intermediate_wire_3[1268]),.o(intermediate_reg_3[634])); 
xor_module xor_module_inst_3_190(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1267]),.i2(intermediate_wire_3[1266]),.o(intermediate_reg_3[633])); 
mux_module mux_module_inst_3_191(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1265]),.i2(intermediate_wire_3[1264]),.o(intermediate_reg_3[632]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_192(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1263]),.i2(intermediate_wire_3[1262]),.o(intermediate_reg_3[631])); 
xor_module xor_module_inst_3_193(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1261]),.i2(intermediate_wire_3[1260]),.o(intermediate_reg_3[630])); 
mux_module mux_module_inst_3_194(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1259]),.i2(intermediate_wire_3[1258]),.o(intermediate_reg_3[629]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_195(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1257]),.i2(intermediate_wire_3[1256]),.o(intermediate_reg_3[628])); 
xor_module xor_module_inst_3_196(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1255]),.i2(intermediate_wire_3[1254]),.o(intermediate_reg_3[627])); 
mux_module mux_module_inst_3_197(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1253]),.i2(intermediate_wire_3[1252]),.o(intermediate_reg_3[626]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_198(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1251]),.i2(intermediate_wire_3[1250]),.o(intermediate_reg_3[625]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_199(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1249]),.i2(intermediate_wire_3[1248]),.o(intermediate_reg_3[624])); 
mux_module mux_module_inst_3_200(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1247]),.i2(intermediate_wire_3[1246]),.o(intermediate_reg_3[623]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_201(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1245]),.i2(intermediate_wire_3[1244]),.o(intermediate_reg_3[622]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_202(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1243]),.i2(intermediate_wire_3[1242]),.o(intermediate_reg_3[621]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_203(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1241]),.i2(intermediate_wire_3[1240]),.o(intermediate_reg_3[620]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_204(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1239]),.i2(intermediate_wire_3[1238]),.o(intermediate_reg_3[619]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_205(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1237]),.i2(intermediate_wire_3[1236]),.o(intermediate_reg_3[618]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_206(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1235]),.i2(intermediate_wire_3[1234]),.o(intermediate_reg_3[617]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_207(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1233]),.i2(intermediate_wire_3[1232]),.o(intermediate_reg_3[616])); 
mux_module mux_module_inst_3_208(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1231]),.i2(intermediate_wire_3[1230]),.o(intermediate_reg_3[615]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_209(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1229]),.i2(intermediate_wire_3[1228]),.o(intermediate_reg_3[614])); 
mux_module mux_module_inst_3_210(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1227]),.i2(intermediate_wire_3[1226]),.o(intermediate_reg_3[613]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_211(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1225]),.i2(intermediate_wire_3[1224]),.o(intermediate_reg_3[612]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_212(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1223]),.i2(intermediate_wire_3[1222]),.o(intermediate_reg_3[611]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_213(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1221]),.i2(intermediate_wire_3[1220]),.o(intermediate_reg_3[610])); 
mux_module mux_module_inst_3_214(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1219]),.i2(intermediate_wire_3[1218]),.o(intermediate_reg_3[609]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_215(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1217]),.i2(intermediate_wire_3[1216]),.o(intermediate_reg_3[608]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_216(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1215]),.i2(intermediate_wire_3[1214]),.o(intermediate_reg_3[607])); 
mux_module mux_module_inst_3_217(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1213]),.i2(intermediate_wire_3[1212]),.o(intermediate_reg_3[606]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_218(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1211]),.i2(intermediate_wire_3[1210]),.o(intermediate_reg_3[605]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_219(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1209]),.i2(intermediate_wire_3[1208]),.o(intermediate_reg_3[604]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_220(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1207]),.i2(intermediate_wire_3[1206]),.o(intermediate_reg_3[603])); 
mux_module mux_module_inst_3_221(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1205]),.i2(intermediate_wire_3[1204]),.o(intermediate_reg_3[602]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_222(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1203]),.i2(intermediate_wire_3[1202]),.o(intermediate_reg_3[601])); 
mux_module mux_module_inst_3_223(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1201]),.i2(intermediate_wire_3[1200]),.o(intermediate_reg_3[600]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_224(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1199]),.i2(intermediate_wire_3[1198]),.o(intermediate_reg_3[599])); 
xor_module xor_module_inst_3_225(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1197]),.i2(intermediate_wire_3[1196]),.o(intermediate_reg_3[598])); 
mux_module mux_module_inst_3_226(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1195]),.i2(intermediate_wire_3[1194]),.o(intermediate_reg_3[597]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_227(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1193]),.i2(intermediate_wire_3[1192]),.o(intermediate_reg_3[596]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_228(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1191]),.i2(intermediate_wire_3[1190]),.o(intermediate_reg_3[595]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_229(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1189]),.i2(intermediate_wire_3[1188]),.o(intermediate_reg_3[594]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_230(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1187]),.i2(intermediate_wire_3[1186]),.o(intermediate_reg_3[593])); 
xor_module xor_module_inst_3_231(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1185]),.i2(intermediate_wire_3[1184]),.o(intermediate_reg_3[592])); 
xor_module xor_module_inst_3_232(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1183]),.i2(intermediate_wire_3[1182]),.o(intermediate_reg_3[591])); 
xor_module xor_module_inst_3_233(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1181]),.i2(intermediate_wire_3[1180]),.o(intermediate_reg_3[590])); 
xor_module xor_module_inst_3_234(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1179]),.i2(intermediate_wire_3[1178]),.o(intermediate_reg_3[589])); 
mux_module mux_module_inst_3_235(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1177]),.i2(intermediate_wire_3[1176]),.o(intermediate_reg_3[588]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_236(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1175]),.i2(intermediate_wire_3[1174]),.o(intermediate_reg_3[587])); 
xor_module xor_module_inst_3_237(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1173]),.i2(intermediate_wire_3[1172]),.o(intermediate_reg_3[586])); 
xor_module xor_module_inst_3_238(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1171]),.i2(intermediate_wire_3[1170]),.o(intermediate_reg_3[585])); 
mux_module mux_module_inst_3_239(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1169]),.i2(intermediate_wire_3[1168]),.o(intermediate_reg_3[584]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_240(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1167]),.i2(intermediate_wire_3[1166]),.o(intermediate_reg_3[583]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_241(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1165]),.i2(intermediate_wire_3[1164]),.o(intermediate_reg_3[582])); 
mux_module mux_module_inst_3_242(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1163]),.i2(intermediate_wire_3[1162]),.o(intermediate_reg_3[581]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_243(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1161]),.i2(intermediate_wire_3[1160]),.o(intermediate_reg_3[580])); 
mux_module mux_module_inst_3_244(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1159]),.i2(intermediate_wire_3[1158]),.o(intermediate_reg_3[579]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_245(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1157]),.i2(intermediate_wire_3[1156]),.o(intermediate_reg_3[578])); 
mux_module mux_module_inst_3_246(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1155]),.i2(intermediate_wire_3[1154]),.o(intermediate_reg_3[577]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_247(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1153]),.i2(intermediate_wire_3[1152]),.o(intermediate_reg_3[576]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_248(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1151]),.i2(intermediate_wire_3[1150]),.o(intermediate_reg_3[575])); 
mux_module mux_module_inst_3_249(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1149]),.i2(intermediate_wire_3[1148]),.o(intermediate_reg_3[574]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_250(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1147]),.i2(intermediate_wire_3[1146]),.o(intermediate_reg_3[573]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_251(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1145]),.i2(intermediate_wire_3[1144]),.o(intermediate_reg_3[572])); 
mux_module mux_module_inst_3_252(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1143]),.i2(intermediate_wire_3[1142]),.o(intermediate_reg_3[571]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_253(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1141]),.i2(intermediate_wire_3[1140]),.o(intermediate_reg_3[570]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_254(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1139]),.i2(intermediate_wire_3[1138]),.o(intermediate_reg_3[569]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_255(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1137]),.i2(intermediate_wire_3[1136]),.o(intermediate_reg_3[568]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_256(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1135]),.i2(intermediate_wire_3[1134]),.o(intermediate_reg_3[567]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_257(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1133]),.i2(intermediate_wire_3[1132]),.o(intermediate_reg_3[566]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_258(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1131]),.i2(intermediate_wire_3[1130]),.o(intermediate_reg_3[565])); 
mux_module mux_module_inst_3_259(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1129]),.i2(intermediate_wire_3[1128]),.o(intermediate_reg_3[564]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_260(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1127]),.i2(intermediate_wire_3[1126]),.o(intermediate_reg_3[563])); 
xor_module xor_module_inst_3_261(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1125]),.i2(intermediate_wire_3[1124]),.o(intermediate_reg_3[562])); 
xor_module xor_module_inst_3_262(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1123]),.i2(intermediate_wire_3[1122]),.o(intermediate_reg_3[561])); 
xor_module xor_module_inst_3_263(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1121]),.i2(intermediate_wire_3[1120]),.o(intermediate_reg_3[560])); 
mux_module mux_module_inst_3_264(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1119]),.i2(intermediate_wire_3[1118]),.o(intermediate_reg_3[559]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_265(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1117]),.i2(intermediate_wire_3[1116]),.o(intermediate_reg_3[558]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_266(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1115]),.i2(intermediate_wire_3[1114]),.o(intermediate_reg_3[557]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_267(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1113]),.i2(intermediate_wire_3[1112]),.o(intermediate_reg_3[556]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_268(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1111]),.i2(intermediate_wire_3[1110]),.o(intermediate_reg_3[555]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_269(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1109]),.i2(intermediate_wire_3[1108]),.o(intermediate_reg_3[554]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_270(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1107]),.i2(intermediate_wire_3[1106]),.o(intermediate_reg_3[553])); 
mux_module mux_module_inst_3_271(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1105]),.i2(intermediate_wire_3[1104]),.o(intermediate_reg_3[552]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_272(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1103]),.i2(intermediate_wire_3[1102]),.o(intermediate_reg_3[551])); 
xor_module xor_module_inst_3_273(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1101]),.i2(intermediate_wire_3[1100]),.o(intermediate_reg_3[550])); 
xor_module xor_module_inst_3_274(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1099]),.i2(intermediate_wire_3[1098]),.o(intermediate_reg_3[549])); 
xor_module xor_module_inst_3_275(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1097]),.i2(intermediate_wire_3[1096]),.o(intermediate_reg_3[548])); 
mux_module mux_module_inst_3_276(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1095]),.i2(intermediate_wire_3[1094]),.o(intermediate_reg_3[547]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_277(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1093]),.i2(intermediate_wire_3[1092]),.o(intermediate_reg_3[546])); 
xor_module xor_module_inst_3_278(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1091]),.i2(intermediate_wire_3[1090]),.o(intermediate_reg_3[545])); 
xor_module xor_module_inst_3_279(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1089]),.i2(intermediate_wire_3[1088]),.o(intermediate_reg_3[544])); 
mux_module mux_module_inst_3_280(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1087]),.i2(intermediate_wire_3[1086]),.o(intermediate_reg_3[543]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_281(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1085]),.i2(intermediate_wire_3[1084]),.o(intermediate_reg_3[542]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_282(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1083]),.i2(intermediate_wire_3[1082]),.o(intermediate_reg_3[541]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_283(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1081]),.i2(intermediate_wire_3[1080]),.o(intermediate_reg_3[540])); 
xor_module xor_module_inst_3_284(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1079]),.i2(intermediate_wire_3[1078]),.o(intermediate_reg_3[539])); 
xor_module xor_module_inst_3_285(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1077]),.i2(intermediate_wire_3[1076]),.o(intermediate_reg_3[538])); 
mux_module mux_module_inst_3_286(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1075]),.i2(intermediate_wire_3[1074]),.o(intermediate_reg_3[537]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_287(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1073]),.i2(intermediate_wire_3[1072]),.o(intermediate_reg_3[536]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_288(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1071]),.i2(intermediate_wire_3[1070]),.o(intermediate_reg_3[535])); 
mux_module mux_module_inst_3_289(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1069]),.i2(intermediate_wire_3[1068]),.o(intermediate_reg_3[534]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_290(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1067]),.i2(intermediate_wire_3[1066]),.o(intermediate_reg_3[533])); 
xor_module xor_module_inst_3_291(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1065]),.i2(intermediate_wire_3[1064]),.o(intermediate_reg_3[532])); 
mux_module mux_module_inst_3_292(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1063]),.i2(intermediate_wire_3[1062]),.o(intermediate_reg_3[531]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_293(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1061]),.i2(intermediate_wire_3[1060]),.o(intermediate_reg_3[530])); 
mux_module mux_module_inst_3_294(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1059]),.i2(intermediate_wire_3[1058]),.o(intermediate_reg_3[529]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_295(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1057]),.i2(intermediate_wire_3[1056]),.o(intermediate_reg_3[528]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_296(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1055]),.i2(intermediate_wire_3[1054]),.o(intermediate_reg_3[527]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_297(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1053]),.i2(intermediate_wire_3[1052]),.o(intermediate_reg_3[526])); 
mux_module mux_module_inst_3_298(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1051]),.i2(intermediate_wire_3[1050]),.o(intermediate_reg_3[525]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_299(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1049]),.i2(intermediate_wire_3[1048]),.o(intermediate_reg_3[524])); 
mux_module mux_module_inst_3_300(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1047]),.i2(intermediate_wire_3[1046]),.o(intermediate_reg_3[523]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_301(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1045]),.i2(intermediate_wire_3[1044]),.o(intermediate_reg_3[522])); 
mux_module mux_module_inst_3_302(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1043]),.i2(intermediate_wire_3[1042]),.o(intermediate_reg_3[521]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_303(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1041]),.i2(intermediate_wire_3[1040]),.o(intermediate_reg_3[520])); 
mux_module mux_module_inst_3_304(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1039]),.i2(intermediate_wire_3[1038]),.o(intermediate_reg_3[519]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_305(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1037]),.i2(intermediate_wire_3[1036]),.o(intermediate_reg_3[518]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_306(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1035]),.i2(intermediate_wire_3[1034]),.o(intermediate_reg_3[517]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_307(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1033]),.i2(intermediate_wire_3[1032]),.o(intermediate_reg_3[516]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_308(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1031]),.i2(intermediate_wire_3[1030]),.o(intermediate_reg_3[515])); 
mux_module mux_module_inst_3_309(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1029]),.i2(intermediate_wire_3[1028]),.o(intermediate_reg_3[514]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_310(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1027]),.i2(intermediate_wire_3[1026]),.o(intermediate_reg_3[513])); 
mux_module mux_module_inst_3_311(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1025]),.i2(intermediate_wire_3[1024]),.o(intermediate_reg_3[512]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_312(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1023]),.i2(intermediate_wire_3[1022]),.o(intermediate_reg_3[511]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_313(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1021]),.i2(intermediate_wire_3[1020]),.o(intermediate_reg_3[510]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_314(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1019]),.i2(intermediate_wire_3[1018]),.o(intermediate_reg_3[509])); 
xor_module xor_module_inst_3_315(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1017]),.i2(intermediate_wire_3[1016]),.o(intermediate_reg_3[508])); 
mux_module mux_module_inst_3_316(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1015]),.i2(intermediate_wire_3[1014]),.o(intermediate_reg_3[507]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_317(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1013]),.i2(intermediate_wire_3[1012]),.o(intermediate_reg_3[506]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_318(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1011]),.i2(intermediate_wire_3[1010]),.o(intermediate_reg_3[505]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_319(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1009]),.i2(intermediate_wire_3[1008]),.o(intermediate_reg_3[504])); 
xor_module xor_module_inst_3_320(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1007]),.i2(intermediate_wire_3[1006]),.o(intermediate_reg_3[503])); 
xor_module xor_module_inst_3_321(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1005]),.i2(intermediate_wire_3[1004]),.o(intermediate_reg_3[502])); 
xor_module xor_module_inst_3_322(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1003]),.i2(intermediate_wire_3[1002]),.o(intermediate_reg_3[501])); 
mux_module mux_module_inst_3_323(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1001]),.i2(intermediate_wire_3[1000]),.o(intermediate_reg_3[500]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_324(.clk(clk),.reset(reset),.i1(intermediate_wire_3[999]),.i2(intermediate_wire_3[998]),.o(intermediate_reg_3[499])); 
mux_module mux_module_inst_3_325(.clk(clk),.reset(reset),.i1(intermediate_wire_3[997]),.i2(intermediate_wire_3[996]),.o(intermediate_reg_3[498]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_326(.clk(clk),.reset(reset),.i1(intermediate_wire_3[995]),.i2(intermediate_wire_3[994]),.o(intermediate_reg_3[497])); 
mux_module mux_module_inst_3_327(.clk(clk),.reset(reset),.i1(intermediate_wire_3[993]),.i2(intermediate_wire_3[992]),.o(intermediate_reg_3[496]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_328(.clk(clk),.reset(reset),.i1(intermediate_wire_3[991]),.i2(intermediate_wire_3[990]),.o(intermediate_reg_3[495]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_329(.clk(clk),.reset(reset),.i1(intermediate_wire_3[989]),.i2(intermediate_wire_3[988]),.o(intermediate_reg_3[494]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_330(.clk(clk),.reset(reset),.i1(intermediate_wire_3[987]),.i2(intermediate_wire_3[986]),.o(intermediate_reg_3[493]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_331(.clk(clk),.reset(reset),.i1(intermediate_wire_3[985]),.i2(intermediate_wire_3[984]),.o(intermediate_reg_3[492]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_332(.clk(clk),.reset(reset),.i1(intermediate_wire_3[983]),.i2(intermediate_wire_3[982]),.o(intermediate_reg_3[491]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_333(.clk(clk),.reset(reset),.i1(intermediate_wire_3[981]),.i2(intermediate_wire_3[980]),.o(intermediate_reg_3[490]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_334(.clk(clk),.reset(reset),.i1(intermediate_wire_3[979]),.i2(intermediate_wire_3[978]),.o(intermediate_reg_3[489]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_335(.clk(clk),.reset(reset),.i1(intermediate_wire_3[977]),.i2(intermediate_wire_3[976]),.o(intermediate_reg_3[488])); 
mux_module mux_module_inst_3_336(.clk(clk),.reset(reset),.i1(intermediate_wire_3[975]),.i2(intermediate_wire_3[974]),.o(intermediate_reg_3[487]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_337(.clk(clk),.reset(reset),.i1(intermediate_wire_3[973]),.i2(intermediate_wire_3[972]),.o(intermediate_reg_3[486])); 
xor_module xor_module_inst_3_338(.clk(clk),.reset(reset),.i1(intermediate_wire_3[971]),.i2(intermediate_wire_3[970]),.o(intermediate_reg_3[485])); 
mux_module mux_module_inst_3_339(.clk(clk),.reset(reset),.i1(intermediate_wire_3[969]),.i2(intermediate_wire_3[968]),.o(intermediate_reg_3[484]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_340(.clk(clk),.reset(reset),.i1(intermediate_wire_3[967]),.i2(intermediate_wire_3[966]),.o(intermediate_reg_3[483]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_341(.clk(clk),.reset(reset),.i1(intermediate_wire_3[965]),.i2(intermediate_wire_3[964]),.o(intermediate_reg_3[482])); 
xor_module xor_module_inst_3_342(.clk(clk),.reset(reset),.i1(intermediate_wire_3[963]),.i2(intermediate_wire_3[962]),.o(intermediate_reg_3[481])); 
xor_module xor_module_inst_3_343(.clk(clk),.reset(reset),.i1(intermediate_wire_3[961]),.i2(intermediate_wire_3[960]),.o(intermediate_reg_3[480])); 
mux_module mux_module_inst_3_344(.clk(clk),.reset(reset),.i1(intermediate_wire_3[959]),.i2(intermediate_wire_3[958]),.o(intermediate_reg_3[479]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_345(.clk(clk),.reset(reset),.i1(intermediate_wire_3[957]),.i2(intermediate_wire_3[956]),.o(intermediate_reg_3[478])); 
xor_module xor_module_inst_3_346(.clk(clk),.reset(reset),.i1(intermediate_wire_3[955]),.i2(intermediate_wire_3[954]),.o(intermediate_reg_3[477])); 
xor_module xor_module_inst_3_347(.clk(clk),.reset(reset),.i1(intermediate_wire_3[953]),.i2(intermediate_wire_3[952]),.o(intermediate_reg_3[476])); 
xor_module xor_module_inst_3_348(.clk(clk),.reset(reset),.i1(intermediate_wire_3[951]),.i2(intermediate_wire_3[950]),.o(intermediate_reg_3[475])); 
mux_module mux_module_inst_3_349(.clk(clk),.reset(reset),.i1(intermediate_wire_3[949]),.i2(intermediate_wire_3[948]),.o(intermediate_reg_3[474]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_350(.clk(clk),.reset(reset),.i1(intermediate_wire_3[947]),.i2(intermediate_wire_3[946]),.o(intermediate_reg_3[473]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_351(.clk(clk),.reset(reset),.i1(intermediate_wire_3[945]),.i2(intermediate_wire_3[944]),.o(intermediate_reg_3[472]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_352(.clk(clk),.reset(reset),.i1(intermediate_wire_3[943]),.i2(intermediate_wire_3[942]),.o(intermediate_reg_3[471])); 
xor_module xor_module_inst_3_353(.clk(clk),.reset(reset),.i1(intermediate_wire_3[941]),.i2(intermediate_wire_3[940]),.o(intermediate_reg_3[470])); 
mux_module mux_module_inst_3_354(.clk(clk),.reset(reset),.i1(intermediate_wire_3[939]),.i2(intermediate_wire_3[938]),.o(intermediate_reg_3[469]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_355(.clk(clk),.reset(reset),.i1(intermediate_wire_3[937]),.i2(intermediate_wire_3[936]),.o(intermediate_reg_3[468])); 
xor_module xor_module_inst_3_356(.clk(clk),.reset(reset),.i1(intermediate_wire_3[935]),.i2(intermediate_wire_3[934]),.o(intermediate_reg_3[467])); 
mux_module mux_module_inst_3_357(.clk(clk),.reset(reset),.i1(intermediate_wire_3[933]),.i2(intermediate_wire_3[932]),.o(intermediate_reg_3[466]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_358(.clk(clk),.reset(reset),.i1(intermediate_wire_3[931]),.i2(intermediate_wire_3[930]),.o(intermediate_reg_3[465])); 
xor_module xor_module_inst_3_359(.clk(clk),.reset(reset),.i1(intermediate_wire_3[929]),.i2(intermediate_wire_3[928]),.o(intermediate_reg_3[464])); 
mux_module mux_module_inst_3_360(.clk(clk),.reset(reset),.i1(intermediate_wire_3[927]),.i2(intermediate_wire_3[926]),.o(intermediate_reg_3[463]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_361(.clk(clk),.reset(reset),.i1(intermediate_wire_3[925]),.i2(intermediate_wire_3[924]),.o(intermediate_reg_3[462])); 
mux_module mux_module_inst_3_362(.clk(clk),.reset(reset),.i1(intermediate_wire_3[923]),.i2(intermediate_wire_3[922]),.o(intermediate_reg_3[461]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_363(.clk(clk),.reset(reset),.i1(intermediate_wire_3[921]),.i2(intermediate_wire_3[920]),.o(intermediate_reg_3[460])); 
xor_module xor_module_inst_3_364(.clk(clk),.reset(reset),.i1(intermediate_wire_3[919]),.i2(intermediate_wire_3[918]),.o(intermediate_reg_3[459])); 
mux_module mux_module_inst_3_365(.clk(clk),.reset(reset),.i1(intermediate_wire_3[917]),.i2(intermediate_wire_3[916]),.o(intermediate_reg_3[458]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_366(.clk(clk),.reset(reset),.i1(intermediate_wire_3[915]),.i2(intermediate_wire_3[914]),.o(intermediate_reg_3[457])); 
mux_module mux_module_inst_3_367(.clk(clk),.reset(reset),.i1(intermediate_wire_3[913]),.i2(intermediate_wire_3[912]),.o(intermediate_reg_3[456]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_368(.clk(clk),.reset(reset),.i1(intermediate_wire_3[911]),.i2(intermediate_wire_3[910]),.o(intermediate_reg_3[455])); 
xor_module xor_module_inst_3_369(.clk(clk),.reset(reset),.i1(intermediate_wire_3[909]),.i2(intermediate_wire_3[908]),.o(intermediate_reg_3[454])); 
mux_module mux_module_inst_3_370(.clk(clk),.reset(reset),.i1(intermediate_wire_3[907]),.i2(intermediate_wire_3[906]),.o(intermediate_reg_3[453]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_371(.clk(clk),.reset(reset),.i1(intermediate_wire_3[905]),.i2(intermediate_wire_3[904]),.o(intermediate_reg_3[452])); 
xor_module xor_module_inst_3_372(.clk(clk),.reset(reset),.i1(intermediate_wire_3[903]),.i2(intermediate_wire_3[902]),.o(intermediate_reg_3[451])); 
xor_module xor_module_inst_3_373(.clk(clk),.reset(reset),.i1(intermediate_wire_3[901]),.i2(intermediate_wire_3[900]),.o(intermediate_reg_3[450])); 
mux_module mux_module_inst_3_374(.clk(clk),.reset(reset),.i1(intermediate_wire_3[899]),.i2(intermediate_wire_3[898]),.o(intermediate_reg_3[449]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_375(.clk(clk),.reset(reset),.i1(intermediate_wire_3[897]),.i2(intermediate_wire_3[896]),.o(intermediate_reg_3[448]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_376(.clk(clk),.reset(reset),.i1(intermediate_wire_3[895]),.i2(intermediate_wire_3[894]),.o(intermediate_reg_3[447]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_377(.clk(clk),.reset(reset),.i1(intermediate_wire_3[893]),.i2(intermediate_wire_3[892]),.o(intermediate_reg_3[446]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_378(.clk(clk),.reset(reset),.i1(intermediate_wire_3[891]),.i2(intermediate_wire_3[890]),.o(intermediate_reg_3[445])); 
mux_module mux_module_inst_3_379(.clk(clk),.reset(reset),.i1(intermediate_wire_3[889]),.i2(intermediate_wire_3[888]),.o(intermediate_reg_3[444]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_380(.clk(clk),.reset(reset),.i1(intermediate_wire_3[887]),.i2(intermediate_wire_3[886]),.o(intermediate_reg_3[443])); 
mux_module mux_module_inst_3_381(.clk(clk),.reset(reset),.i1(intermediate_wire_3[885]),.i2(intermediate_wire_3[884]),.o(intermediate_reg_3[442]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_382(.clk(clk),.reset(reset),.i1(intermediate_wire_3[883]),.i2(intermediate_wire_3[882]),.o(intermediate_reg_3[441]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_383(.clk(clk),.reset(reset),.i1(intermediate_wire_3[881]),.i2(intermediate_wire_3[880]),.o(intermediate_reg_3[440]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_384(.clk(clk),.reset(reset),.i1(intermediate_wire_3[879]),.i2(intermediate_wire_3[878]),.o(intermediate_reg_3[439]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_385(.clk(clk),.reset(reset),.i1(intermediate_wire_3[877]),.i2(intermediate_wire_3[876]),.o(intermediate_reg_3[438])); 
xor_module xor_module_inst_3_386(.clk(clk),.reset(reset),.i1(intermediate_wire_3[875]),.i2(intermediate_wire_3[874]),.o(intermediate_reg_3[437])); 
xor_module xor_module_inst_3_387(.clk(clk),.reset(reset),.i1(intermediate_wire_3[873]),.i2(intermediate_wire_3[872]),.o(intermediate_reg_3[436])); 
xor_module xor_module_inst_3_388(.clk(clk),.reset(reset),.i1(intermediate_wire_3[871]),.i2(intermediate_wire_3[870]),.o(intermediate_reg_3[435])); 
xor_module xor_module_inst_3_389(.clk(clk),.reset(reset),.i1(intermediate_wire_3[869]),.i2(intermediate_wire_3[868]),.o(intermediate_reg_3[434])); 
mux_module mux_module_inst_3_390(.clk(clk),.reset(reset),.i1(intermediate_wire_3[867]),.i2(intermediate_wire_3[866]),.o(intermediate_reg_3[433]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_391(.clk(clk),.reset(reset),.i1(intermediate_wire_3[865]),.i2(intermediate_wire_3[864]),.o(intermediate_reg_3[432]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_392(.clk(clk),.reset(reset),.i1(intermediate_wire_3[863]),.i2(intermediate_wire_3[862]),.o(intermediate_reg_3[431]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_393(.clk(clk),.reset(reset),.i1(intermediate_wire_3[861]),.i2(intermediate_wire_3[860]),.o(intermediate_reg_3[430]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_394(.clk(clk),.reset(reset),.i1(intermediate_wire_3[859]),.i2(intermediate_wire_3[858]),.o(intermediate_reg_3[429])); 
mux_module mux_module_inst_3_395(.clk(clk),.reset(reset),.i1(intermediate_wire_3[857]),.i2(intermediate_wire_3[856]),.o(intermediate_reg_3[428]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_396(.clk(clk),.reset(reset),.i1(intermediate_wire_3[855]),.i2(intermediate_wire_3[854]),.o(intermediate_reg_3[427]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_397(.clk(clk),.reset(reset),.i1(intermediate_wire_3[853]),.i2(intermediate_wire_3[852]),.o(intermediate_reg_3[426])); 
mux_module mux_module_inst_3_398(.clk(clk),.reset(reset),.i1(intermediate_wire_3[851]),.i2(intermediate_wire_3[850]),.o(intermediate_reg_3[425]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_399(.clk(clk),.reset(reset),.i1(intermediate_wire_3[849]),.i2(intermediate_wire_3[848]),.o(intermediate_reg_3[424])); 
xor_module xor_module_inst_3_400(.clk(clk),.reset(reset),.i1(intermediate_wire_3[847]),.i2(intermediate_wire_3[846]),.o(intermediate_reg_3[423])); 
xor_module xor_module_inst_3_401(.clk(clk),.reset(reset),.i1(intermediate_wire_3[845]),.i2(intermediate_wire_3[844]),.o(intermediate_reg_3[422])); 
xor_module xor_module_inst_3_402(.clk(clk),.reset(reset),.i1(intermediate_wire_3[843]),.i2(intermediate_wire_3[842]),.o(intermediate_reg_3[421])); 
xor_module xor_module_inst_3_403(.clk(clk),.reset(reset),.i1(intermediate_wire_3[841]),.i2(intermediate_wire_3[840]),.o(intermediate_reg_3[420])); 
xor_module xor_module_inst_3_404(.clk(clk),.reset(reset),.i1(intermediate_wire_3[839]),.i2(intermediate_wire_3[838]),.o(intermediate_reg_3[419])); 
xor_module xor_module_inst_3_405(.clk(clk),.reset(reset),.i1(intermediate_wire_3[837]),.i2(intermediate_wire_3[836]),.o(intermediate_reg_3[418])); 
xor_module xor_module_inst_3_406(.clk(clk),.reset(reset),.i1(intermediate_wire_3[835]),.i2(intermediate_wire_3[834]),.o(intermediate_reg_3[417])); 
mux_module mux_module_inst_3_407(.clk(clk),.reset(reset),.i1(intermediate_wire_3[833]),.i2(intermediate_wire_3[832]),.o(intermediate_reg_3[416]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_408(.clk(clk),.reset(reset),.i1(intermediate_wire_3[831]),.i2(intermediate_wire_3[830]),.o(intermediate_reg_3[415]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_409(.clk(clk),.reset(reset),.i1(intermediate_wire_3[829]),.i2(intermediate_wire_3[828]),.o(intermediate_reg_3[414]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_410(.clk(clk),.reset(reset),.i1(intermediate_wire_3[827]),.i2(intermediate_wire_3[826]),.o(intermediate_reg_3[413])); 
xor_module xor_module_inst_3_411(.clk(clk),.reset(reset),.i1(intermediate_wire_3[825]),.i2(intermediate_wire_3[824]),.o(intermediate_reg_3[412])); 
xor_module xor_module_inst_3_412(.clk(clk),.reset(reset),.i1(intermediate_wire_3[823]),.i2(intermediate_wire_3[822]),.o(intermediate_reg_3[411])); 
xor_module xor_module_inst_3_413(.clk(clk),.reset(reset),.i1(intermediate_wire_3[821]),.i2(intermediate_wire_3[820]),.o(intermediate_reg_3[410])); 
xor_module xor_module_inst_3_414(.clk(clk),.reset(reset),.i1(intermediate_wire_3[819]),.i2(intermediate_wire_3[818]),.o(intermediate_reg_3[409])); 
xor_module xor_module_inst_3_415(.clk(clk),.reset(reset),.i1(intermediate_wire_3[817]),.i2(intermediate_wire_3[816]),.o(intermediate_reg_3[408])); 
mux_module mux_module_inst_3_416(.clk(clk),.reset(reset),.i1(intermediate_wire_3[815]),.i2(intermediate_wire_3[814]),.o(intermediate_reg_3[407]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_417(.clk(clk),.reset(reset),.i1(intermediate_wire_3[813]),.i2(intermediate_wire_3[812]),.o(intermediate_reg_3[406])); 
mux_module mux_module_inst_3_418(.clk(clk),.reset(reset),.i1(intermediate_wire_3[811]),.i2(intermediate_wire_3[810]),.o(intermediate_reg_3[405]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_419(.clk(clk),.reset(reset),.i1(intermediate_wire_3[809]),.i2(intermediate_wire_3[808]),.o(intermediate_reg_3[404])); 
xor_module xor_module_inst_3_420(.clk(clk),.reset(reset),.i1(intermediate_wire_3[807]),.i2(intermediate_wire_3[806]),.o(intermediate_reg_3[403])); 
mux_module mux_module_inst_3_421(.clk(clk),.reset(reset),.i1(intermediate_wire_3[805]),.i2(intermediate_wire_3[804]),.o(intermediate_reg_3[402]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_422(.clk(clk),.reset(reset),.i1(intermediate_wire_3[803]),.i2(intermediate_wire_3[802]),.o(intermediate_reg_3[401])); 
mux_module mux_module_inst_3_423(.clk(clk),.reset(reset),.i1(intermediate_wire_3[801]),.i2(intermediate_wire_3[800]),.o(intermediate_reg_3[400]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_424(.clk(clk),.reset(reset),.i1(intermediate_wire_3[799]),.i2(intermediate_wire_3[798]),.o(intermediate_reg_3[399]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_425(.clk(clk),.reset(reset),.i1(intermediate_wire_3[797]),.i2(intermediate_wire_3[796]),.o(intermediate_reg_3[398]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_426(.clk(clk),.reset(reset),.i1(intermediate_wire_3[795]),.i2(intermediate_wire_3[794]),.o(intermediate_reg_3[397]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_427(.clk(clk),.reset(reset),.i1(intermediate_wire_3[793]),.i2(intermediate_wire_3[792]),.o(intermediate_reg_3[396]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_428(.clk(clk),.reset(reset),.i1(intermediate_wire_3[791]),.i2(intermediate_wire_3[790]),.o(intermediate_reg_3[395]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_429(.clk(clk),.reset(reset),.i1(intermediate_wire_3[789]),.i2(intermediate_wire_3[788]),.o(intermediate_reg_3[394]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_430(.clk(clk),.reset(reset),.i1(intermediate_wire_3[787]),.i2(intermediate_wire_3[786]),.o(intermediate_reg_3[393]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_431(.clk(clk),.reset(reset),.i1(intermediate_wire_3[785]),.i2(intermediate_wire_3[784]),.o(intermediate_reg_3[392]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_432(.clk(clk),.reset(reset),.i1(intermediate_wire_3[783]),.i2(intermediate_wire_3[782]),.o(intermediate_reg_3[391])); 
xor_module xor_module_inst_3_433(.clk(clk),.reset(reset),.i1(intermediate_wire_3[781]),.i2(intermediate_wire_3[780]),.o(intermediate_reg_3[390])); 
mux_module mux_module_inst_3_434(.clk(clk),.reset(reset),.i1(intermediate_wire_3[779]),.i2(intermediate_wire_3[778]),.o(intermediate_reg_3[389]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_435(.clk(clk),.reset(reset),.i1(intermediate_wire_3[777]),.i2(intermediate_wire_3[776]),.o(intermediate_reg_3[388])); 
xor_module xor_module_inst_3_436(.clk(clk),.reset(reset),.i1(intermediate_wire_3[775]),.i2(intermediate_wire_3[774]),.o(intermediate_reg_3[387])); 
mux_module mux_module_inst_3_437(.clk(clk),.reset(reset),.i1(intermediate_wire_3[773]),.i2(intermediate_wire_3[772]),.o(intermediate_reg_3[386]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_438(.clk(clk),.reset(reset),.i1(intermediate_wire_3[771]),.i2(intermediate_wire_3[770]),.o(intermediate_reg_3[385]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_439(.clk(clk),.reset(reset),.i1(intermediate_wire_3[769]),.i2(intermediate_wire_3[768]),.o(intermediate_reg_3[384])); 
mux_module mux_module_inst_3_440(.clk(clk),.reset(reset),.i1(intermediate_wire_3[767]),.i2(intermediate_wire_3[766]),.o(intermediate_reg_3[383]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_441(.clk(clk),.reset(reset),.i1(intermediate_wire_3[765]),.i2(intermediate_wire_3[764]),.o(intermediate_reg_3[382])); 
xor_module xor_module_inst_3_442(.clk(clk),.reset(reset),.i1(intermediate_wire_3[763]),.i2(intermediate_wire_3[762]),.o(intermediate_reg_3[381])); 
mux_module mux_module_inst_3_443(.clk(clk),.reset(reset),.i1(intermediate_wire_3[761]),.i2(intermediate_wire_3[760]),.o(intermediate_reg_3[380]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_444(.clk(clk),.reset(reset),.i1(intermediate_wire_3[759]),.i2(intermediate_wire_3[758]),.o(intermediate_reg_3[379]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_445(.clk(clk),.reset(reset),.i1(intermediate_wire_3[757]),.i2(intermediate_wire_3[756]),.o(intermediate_reg_3[378]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_446(.clk(clk),.reset(reset),.i1(intermediate_wire_3[755]),.i2(intermediate_wire_3[754]),.o(intermediate_reg_3[377]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_447(.clk(clk),.reset(reset),.i1(intermediate_wire_3[753]),.i2(intermediate_wire_3[752]),.o(intermediate_reg_3[376]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_448(.clk(clk),.reset(reset),.i1(intermediate_wire_3[751]),.i2(intermediate_wire_3[750]),.o(intermediate_reg_3[375])); 
mux_module mux_module_inst_3_449(.clk(clk),.reset(reset),.i1(intermediate_wire_3[749]),.i2(intermediate_wire_3[748]),.o(intermediate_reg_3[374]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_450(.clk(clk),.reset(reset),.i1(intermediate_wire_3[747]),.i2(intermediate_wire_3[746]),.o(intermediate_reg_3[373]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_451(.clk(clk),.reset(reset),.i1(intermediate_wire_3[745]),.i2(intermediate_wire_3[744]),.o(intermediate_reg_3[372]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_452(.clk(clk),.reset(reset),.i1(intermediate_wire_3[743]),.i2(intermediate_wire_3[742]),.o(intermediate_reg_3[371]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_453(.clk(clk),.reset(reset),.i1(intermediate_wire_3[741]),.i2(intermediate_wire_3[740]),.o(intermediate_reg_3[370])); 
xor_module xor_module_inst_3_454(.clk(clk),.reset(reset),.i1(intermediate_wire_3[739]),.i2(intermediate_wire_3[738]),.o(intermediate_reg_3[369])); 
xor_module xor_module_inst_3_455(.clk(clk),.reset(reset),.i1(intermediate_wire_3[737]),.i2(intermediate_wire_3[736]),.o(intermediate_reg_3[368])); 
xor_module xor_module_inst_3_456(.clk(clk),.reset(reset),.i1(intermediate_wire_3[735]),.i2(intermediate_wire_3[734]),.o(intermediate_reg_3[367])); 
xor_module xor_module_inst_3_457(.clk(clk),.reset(reset),.i1(intermediate_wire_3[733]),.i2(intermediate_wire_3[732]),.o(intermediate_reg_3[366])); 
xor_module xor_module_inst_3_458(.clk(clk),.reset(reset),.i1(intermediate_wire_3[731]),.i2(intermediate_wire_3[730]),.o(intermediate_reg_3[365])); 
xor_module xor_module_inst_3_459(.clk(clk),.reset(reset),.i1(intermediate_wire_3[729]),.i2(intermediate_wire_3[728]),.o(intermediate_reg_3[364])); 
xor_module xor_module_inst_3_460(.clk(clk),.reset(reset),.i1(intermediate_wire_3[727]),.i2(intermediate_wire_3[726]),.o(intermediate_reg_3[363])); 
mux_module mux_module_inst_3_461(.clk(clk),.reset(reset),.i1(intermediate_wire_3[725]),.i2(intermediate_wire_3[724]),.o(intermediate_reg_3[362]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_462(.clk(clk),.reset(reset),.i1(intermediate_wire_3[723]),.i2(intermediate_wire_3[722]),.o(intermediate_reg_3[361])); 
xor_module xor_module_inst_3_463(.clk(clk),.reset(reset),.i1(intermediate_wire_3[721]),.i2(intermediate_wire_3[720]),.o(intermediate_reg_3[360])); 
xor_module xor_module_inst_3_464(.clk(clk),.reset(reset),.i1(intermediate_wire_3[719]),.i2(intermediate_wire_3[718]),.o(intermediate_reg_3[359])); 
mux_module mux_module_inst_3_465(.clk(clk),.reset(reset),.i1(intermediate_wire_3[717]),.i2(intermediate_wire_3[716]),.o(intermediate_reg_3[358]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_466(.clk(clk),.reset(reset),.i1(intermediate_wire_3[715]),.i2(intermediate_wire_3[714]),.o(intermediate_reg_3[357])); 
mux_module mux_module_inst_3_467(.clk(clk),.reset(reset),.i1(intermediate_wire_3[713]),.i2(intermediate_wire_3[712]),.o(intermediate_reg_3[356]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_468(.clk(clk),.reset(reset),.i1(intermediate_wire_3[711]),.i2(intermediate_wire_3[710]),.o(intermediate_reg_3[355])); 
mux_module mux_module_inst_3_469(.clk(clk),.reset(reset),.i1(intermediate_wire_3[709]),.i2(intermediate_wire_3[708]),.o(intermediate_reg_3[354]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_470(.clk(clk),.reset(reset),.i1(intermediate_wire_3[707]),.i2(intermediate_wire_3[706]),.o(intermediate_reg_3[353]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_471(.clk(clk),.reset(reset),.i1(intermediate_wire_3[705]),.i2(intermediate_wire_3[704]),.o(intermediate_reg_3[352])); 
mux_module mux_module_inst_3_472(.clk(clk),.reset(reset),.i1(intermediate_wire_3[703]),.i2(intermediate_wire_3[702]),.o(intermediate_reg_3[351]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_473(.clk(clk),.reset(reset),.i1(intermediate_wire_3[701]),.i2(intermediate_wire_3[700]),.o(intermediate_reg_3[350]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_474(.clk(clk),.reset(reset),.i1(intermediate_wire_3[699]),.i2(intermediate_wire_3[698]),.o(intermediate_reg_3[349]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_475(.clk(clk),.reset(reset),.i1(intermediate_wire_3[697]),.i2(intermediate_wire_3[696]),.o(intermediate_reg_3[348])); 
xor_module xor_module_inst_3_476(.clk(clk),.reset(reset),.i1(intermediate_wire_3[695]),.i2(intermediate_wire_3[694]),.o(intermediate_reg_3[347])); 
mux_module mux_module_inst_3_477(.clk(clk),.reset(reset),.i1(intermediate_wire_3[693]),.i2(intermediate_wire_3[692]),.o(intermediate_reg_3[346]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_478(.clk(clk),.reset(reset),.i1(intermediate_wire_3[691]),.i2(intermediate_wire_3[690]),.o(intermediate_reg_3[345])); 
xor_module xor_module_inst_3_479(.clk(clk),.reset(reset),.i1(intermediate_wire_3[689]),.i2(intermediate_wire_3[688]),.o(intermediate_reg_3[344])); 
mux_module mux_module_inst_3_480(.clk(clk),.reset(reset),.i1(intermediate_wire_3[687]),.i2(intermediate_wire_3[686]),.o(intermediate_reg_3[343]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_481(.clk(clk),.reset(reset),.i1(intermediate_wire_3[685]),.i2(intermediate_wire_3[684]),.o(intermediate_reg_3[342]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_482(.clk(clk),.reset(reset),.i1(intermediate_wire_3[683]),.i2(intermediate_wire_3[682]),.o(intermediate_reg_3[341]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_483(.clk(clk),.reset(reset),.i1(intermediate_wire_3[681]),.i2(intermediate_wire_3[680]),.o(intermediate_reg_3[340])); 
mux_module mux_module_inst_3_484(.clk(clk),.reset(reset),.i1(intermediate_wire_3[679]),.i2(intermediate_wire_3[678]),.o(intermediate_reg_3[339]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_485(.clk(clk),.reset(reset),.i1(intermediate_wire_3[677]),.i2(intermediate_wire_3[676]),.o(intermediate_reg_3[338])); 
xor_module xor_module_inst_3_486(.clk(clk),.reset(reset),.i1(intermediate_wire_3[675]),.i2(intermediate_wire_3[674]),.o(intermediate_reg_3[337])); 
mux_module mux_module_inst_3_487(.clk(clk),.reset(reset),.i1(intermediate_wire_3[673]),.i2(intermediate_wire_3[672]),.o(intermediate_reg_3[336]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_488(.clk(clk),.reset(reset),.i1(intermediate_wire_3[671]),.i2(intermediate_wire_3[670]),.o(intermediate_reg_3[335]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_489(.clk(clk),.reset(reset),.i1(intermediate_wire_3[669]),.i2(intermediate_wire_3[668]),.o(intermediate_reg_3[334]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_490(.clk(clk),.reset(reset),.i1(intermediate_wire_3[667]),.i2(intermediate_wire_3[666]),.o(intermediate_reg_3[333])); 
mux_module mux_module_inst_3_491(.clk(clk),.reset(reset),.i1(intermediate_wire_3[665]),.i2(intermediate_wire_3[664]),.o(intermediate_reg_3[332]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_492(.clk(clk),.reset(reset),.i1(intermediate_wire_3[663]),.i2(intermediate_wire_3[662]),.o(intermediate_reg_3[331])); 
mux_module mux_module_inst_3_493(.clk(clk),.reset(reset),.i1(intermediate_wire_3[661]),.i2(intermediate_wire_3[660]),.o(intermediate_reg_3[330]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_494(.clk(clk),.reset(reset),.i1(intermediate_wire_3[659]),.i2(intermediate_wire_3[658]),.o(intermediate_reg_3[329])); 
xor_module xor_module_inst_3_495(.clk(clk),.reset(reset),.i1(intermediate_wire_3[657]),.i2(intermediate_wire_3[656]),.o(intermediate_reg_3[328])); 
mux_module mux_module_inst_3_496(.clk(clk),.reset(reset),.i1(intermediate_wire_3[655]),.i2(intermediate_wire_3[654]),.o(intermediate_reg_3[327]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_497(.clk(clk),.reset(reset),.i1(intermediate_wire_3[653]),.i2(intermediate_wire_3[652]),.o(intermediate_reg_3[326])); 
mux_module mux_module_inst_3_498(.clk(clk),.reset(reset),.i1(intermediate_wire_3[651]),.i2(intermediate_wire_3[650]),.o(intermediate_reg_3[325]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_499(.clk(clk),.reset(reset),.i1(intermediate_wire_3[649]),.i2(intermediate_wire_3[648]),.o(intermediate_reg_3[324])); 
mux_module mux_module_inst_3_500(.clk(clk),.reset(reset),.i1(intermediate_wire_3[647]),.i2(intermediate_wire_3[646]),.o(intermediate_reg_3[323]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_501(.clk(clk),.reset(reset),.i1(intermediate_wire_3[645]),.i2(intermediate_wire_3[644]),.o(intermediate_reg_3[322]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_502(.clk(clk),.reset(reset),.i1(intermediate_wire_3[643]),.i2(intermediate_wire_3[642]),.o(intermediate_reg_3[321]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_503(.clk(clk),.reset(reset),.i1(intermediate_wire_3[641]),.i2(intermediate_wire_3[640]),.o(intermediate_reg_3[320])); 
mux_module mux_module_inst_3_504(.clk(clk),.reset(reset),.i1(intermediate_wire_3[639]),.i2(intermediate_wire_3[638]),.o(intermediate_reg_3[319]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_505(.clk(clk),.reset(reset),.i1(intermediate_wire_3[637]),.i2(intermediate_wire_3[636]),.o(intermediate_reg_3[318])); 
mux_module mux_module_inst_3_506(.clk(clk),.reset(reset),.i1(intermediate_wire_3[635]),.i2(intermediate_wire_3[634]),.o(intermediate_reg_3[317]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_507(.clk(clk),.reset(reset),.i1(intermediate_wire_3[633]),.i2(intermediate_wire_3[632]),.o(intermediate_reg_3[316]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_508(.clk(clk),.reset(reset),.i1(intermediate_wire_3[631]),.i2(intermediate_wire_3[630]),.o(intermediate_reg_3[315])); 
mux_module mux_module_inst_3_509(.clk(clk),.reset(reset),.i1(intermediate_wire_3[629]),.i2(intermediate_wire_3[628]),.o(intermediate_reg_3[314]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_510(.clk(clk),.reset(reset),.i1(intermediate_wire_3[627]),.i2(intermediate_wire_3[626]),.o(intermediate_reg_3[313])); 
mux_module mux_module_inst_3_511(.clk(clk),.reset(reset),.i1(intermediate_wire_3[625]),.i2(intermediate_wire_3[624]),.o(intermediate_reg_3[312]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_512(.clk(clk),.reset(reset),.i1(intermediate_wire_3[623]),.i2(intermediate_wire_3[622]),.o(intermediate_reg_3[311]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_513(.clk(clk),.reset(reset),.i1(intermediate_wire_3[621]),.i2(intermediate_wire_3[620]),.o(intermediate_reg_3[310])); 
mux_module mux_module_inst_3_514(.clk(clk),.reset(reset),.i1(intermediate_wire_3[619]),.i2(intermediate_wire_3[618]),.o(intermediate_reg_3[309]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_515(.clk(clk),.reset(reset),.i1(intermediate_wire_3[617]),.i2(intermediate_wire_3[616]),.o(intermediate_reg_3[308])); 
xor_module xor_module_inst_3_516(.clk(clk),.reset(reset),.i1(intermediate_wire_3[615]),.i2(intermediate_wire_3[614]),.o(intermediate_reg_3[307])); 
xor_module xor_module_inst_3_517(.clk(clk),.reset(reset),.i1(intermediate_wire_3[613]),.i2(intermediate_wire_3[612]),.o(intermediate_reg_3[306])); 
xor_module xor_module_inst_3_518(.clk(clk),.reset(reset),.i1(intermediate_wire_3[611]),.i2(intermediate_wire_3[610]),.o(intermediate_reg_3[305])); 
xor_module xor_module_inst_3_519(.clk(clk),.reset(reset),.i1(intermediate_wire_3[609]),.i2(intermediate_wire_3[608]),.o(intermediate_reg_3[304])); 
mux_module mux_module_inst_3_520(.clk(clk),.reset(reset),.i1(intermediate_wire_3[607]),.i2(intermediate_wire_3[606]),.o(intermediate_reg_3[303]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_521(.clk(clk),.reset(reset),.i1(intermediate_wire_3[605]),.i2(intermediate_wire_3[604]),.o(intermediate_reg_3[302])); 
mux_module mux_module_inst_3_522(.clk(clk),.reset(reset),.i1(intermediate_wire_3[603]),.i2(intermediate_wire_3[602]),.o(intermediate_reg_3[301]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_523(.clk(clk),.reset(reset),.i1(intermediate_wire_3[601]),.i2(intermediate_wire_3[600]),.o(intermediate_reg_3[300]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_524(.clk(clk),.reset(reset),.i1(intermediate_wire_3[599]),.i2(intermediate_wire_3[598]),.o(intermediate_reg_3[299]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_525(.clk(clk),.reset(reset),.i1(intermediate_wire_3[597]),.i2(intermediate_wire_3[596]),.o(intermediate_reg_3[298]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_526(.clk(clk),.reset(reset),.i1(intermediate_wire_3[595]),.i2(intermediate_wire_3[594]),.o(intermediate_reg_3[297])); 
xor_module xor_module_inst_3_527(.clk(clk),.reset(reset),.i1(intermediate_wire_3[593]),.i2(intermediate_wire_3[592]),.o(intermediate_reg_3[296])); 
mux_module mux_module_inst_3_528(.clk(clk),.reset(reset),.i1(intermediate_wire_3[591]),.i2(intermediate_wire_3[590]),.o(intermediate_reg_3[295]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_529(.clk(clk),.reset(reset),.i1(intermediate_wire_3[589]),.i2(intermediate_wire_3[588]),.o(intermediate_reg_3[294])); 
xor_module xor_module_inst_3_530(.clk(clk),.reset(reset),.i1(intermediate_wire_3[587]),.i2(intermediate_wire_3[586]),.o(intermediate_reg_3[293])); 
mux_module mux_module_inst_3_531(.clk(clk),.reset(reset),.i1(intermediate_wire_3[585]),.i2(intermediate_wire_3[584]),.o(intermediate_reg_3[292]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_532(.clk(clk),.reset(reset),.i1(intermediate_wire_3[583]),.i2(intermediate_wire_3[582]),.o(intermediate_reg_3[291]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_533(.clk(clk),.reset(reset),.i1(intermediate_wire_3[581]),.i2(intermediate_wire_3[580]),.o(intermediate_reg_3[290])); 
mux_module mux_module_inst_3_534(.clk(clk),.reset(reset),.i1(intermediate_wire_3[579]),.i2(intermediate_wire_3[578]),.o(intermediate_reg_3[289]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_535(.clk(clk),.reset(reset),.i1(intermediate_wire_3[577]),.i2(intermediate_wire_3[576]),.o(intermediate_reg_3[288])); 
mux_module mux_module_inst_3_536(.clk(clk),.reset(reset),.i1(intermediate_wire_3[575]),.i2(intermediate_wire_3[574]),.o(intermediate_reg_3[287]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_537(.clk(clk),.reset(reset),.i1(intermediate_wire_3[573]),.i2(intermediate_wire_3[572]),.o(intermediate_reg_3[286]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_538(.clk(clk),.reset(reset),.i1(intermediate_wire_3[571]),.i2(intermediate_wire_3[570]),.o(intermediate_reg_3[285]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_539(.clk(clk),.reset(reset),.i1(intermediate_wire_3[569]),.i2(intermediate_wire_3[568]),.o(intermediate_reg_3[284])); 
xor_module xor_module_inst_3_540(.clk(clk),.reset(reset),.i1(intermediate_wire_3[567]),.i2(intermediate_wire_3[566]),.o(intermediate_reg_3[283])); 
xor_module xor_module_inst_3_541(.clk(clk),.reset(reset),.i1(intermediate_wire_3[565]),.i2(intermediate_wire_3[564]),.o(intermediate_reg_3[282])); 
mux_module mux_module_inst_3_542(.clk(clk),.reset(reset),.i1(intermediate_wire_3[563]),.i2(intermediate_wire_3[562]),.o(intermediate_reg_3[281]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_543(.clk(clk),.reset(reset),.i1(intermediate_wire_3[561]),.i2(intermediate_wire_3[560]),.o(intermediate_reg_3[280]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_544(.clk(clk),.reset(reset),.i1(intermediate_wire_3[559]),.i2(intermediate_wire_3[558]),.o(intermediate_reg_3[279])); 
mux_module mux_module_inst_3_545(.clk(clk),.reset(reset),.i1(intermediate_wire_3[557]),.i2(intermediate_wire_3[556]),.o(intermediate_reg_3[278]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_546(.clk(clk),.reset(reset),.i1(intermediate_wire_3[555]),.i2(intermediate_wire_3[554]),.o(intermediate_reg_3[277])); 
mux_module mux_module_inst_3_547(.clk(clk),.reset(reset),.i1(intermediate_wire_3[553]),.i2(intermediate_wire_3[552]),.o(intermediate_reg_3[276]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_548(.clk(clk),.reset(reset),.i1(intermediate_wire_3[551]),.i2(intermediate_wire_3[550]),.o(intermediate_reg_3[275])); 
mux_module mux_module_inst_3_549(.clk(clk),.reset(reset),.i1(intermediate_wire_3[549]),.i2(intermediate_wire_3[548]),.o(intermediate_reg_3[274]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_550(.clk(clk),.reset(reset),.i1(intermediate_wire_3[547]),.i2(intermediate_wire_3[546]),.o(intermediate_reg_3[273])); 
mux_module mux_module_inst_3_551(.clk(clk),.reset(reset),.i1(intermediate_wire_3[545]),.i2(intermediate_wire_3[544]),.o(intermediate_reg_3[272]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_552(.clk(clk),.reset(reset),.i1(intermediate_wire_3[543]),.i2(intermediate_wire_3[542]),.o(intermediate_reg_3[271])); 
xor_module xor_module_inst_3_553(.clk(clk),.reset(reset),.i1(intermediate_wire_3[541]),.i2(intermediate_wire_3[540]),.o(intermediate_reg_3[270])); 
mux_module mux_module_inst_3_554(.clk(clk),.reset(reset),.i1(intermediate_wire_3[539]),.i2(intermediate_wire_3[538]),.o(intermediate_reg_3[269]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_555(.clk(clk),.reset(reset),.i1(intermediate_wire_3[537]),.i2(intermediate_wire_3[536]),.o(intermediate_reg_3[268])); 
mux_module mux_module_inst_3_556(.clk(clk),.reset(reset),.i1(intermediate_wire_3[535]),.i2(intermediate_wire_3[534]),.o(intermediate_reg_3[267]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_557(.clk(clk),.reset(reset),.i1(intermediate_wire_3[533]),.i2(intermediate_wire_3[532]),.o(intermediate_reg_3[266])); 
xor_module xor_module_inst_3_558(.clk(clk),.reset(reset),.i1(intermediate_wire_3[531]),.i2(intermediate_wire_3[530]),.o(intermediate_reg_3[265])); 
mux_module mux_module_inst_3_559(.clk(clk),.reset(reset),.i1(intermediate_wire_3[529]),.i2(intermediate_wire_3[528]),.o(intermediate_reg_3[264]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_560(.clk(clk),.reset(reset),.i1(intermediate_wire_3[527]),.i2(intermediate_wire_3[526]),.o(intermediate_reg_3[263]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_561(.clk(clk),.reset(reset),.i1(intermediate_wire_3[525]),.i2(intermediate_wire_3[524]),.o(intermediate_reg_3[262])); 
xor_module xor_module_inst_3_562(.clk(clk),.reset(reset),.i1(intermediate_wire_3[523]),.i2(intermediate_wire_3[522]),.o(intermediate_reg_3[261])); 
mux_module mux_module_inst_3_563(.clk(clk),.reset(reset),.i1(intermediate_wire_3[521]),.i2(intermediate_wire_3[520]),.o(intermediate_reg_3[260]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_564(.clk(clk),.reset(reset),.i1(intermediate_wire_3[519]),.i2(intermediate_wire_3[518]),.o(intermediate_reg_3[259])); 
mux_module mux_module_inst_3_565(.clk(clk),.reset(reset),.i1(intermediate_wire_3[517]),.i2(intermediate_wire_3[516]),.o(intermediate_reg_3[258]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_566(.clk(clk),.reset(reset),.i1(intermediate_wire_3[515]),.i2(intermediate_wire_3[514]),.o(intermediate_reg_3[257])); 
mux_module mux_module_inst_3_567(.clk(clk),.reset(reset),.i1(intermediate_wire_3[513]),.i2(intermediate_wire_3[512]),.o(intermediate_reg_3[256]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_568(.clk(clk),.reset(reset),.i1(intermediate_wire_3[511]),.i2(intermediate_wire_3[510]),.o(intermediate_reg_3[255]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_569(.clk(clk),.reset(reset),.i1(intermediate_wire_3[509]),.i2(intermediate_wire_3[508]),.o(intermediate_reg_3[254]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_570(.clk(clk),.reset(reset),.i1(intermediate_wire_3[507]),.i2(intermediate_wire_3[506]),.o(intermediate_reg_3[253])); 
xor_module xor_module_inst_3_571(.clk(clk),.reset(reset),.i1(intermediate_wire_3[505]),.i2(intermediate_wire_3[504]),.o(intermediate_reg_3[252])); 
mux_module mux_module_inst_3_572(.clk(clk),.reset(reset),.i1(intermediate_wire_3[503]),.i2(intermediate_wire_3[502]),.o(intermediate_reg_3[251]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_573(.clk(clk),.reset(reset),.i1(intermediate_wire_3[501]),.i2(intermediate_wire_3[500]),.o(intermediate_reg_3[250]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_574(.clk(clk),.reset(reset),.i1(intermediate_wire_3[499]),.i2(intermediate_wire_3[498]),.o(intermediate_reg_3[249])); 
mux_module mux_module_inst_3_575(.clk(clk),.reset(reset),.i1(intermediate_wire_3[497]),.i2(intermediate_wire_3[496]),.o(intermediate_reg_3[248]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_576(.clk(clk),.reset(reset),.i1(intermediate_wire_3[495]),.i2(intermediate_wire_3[494]),.o(intermediate_reg_3[247]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_577(.clk(clk),.reset(reset),.i1(intermediate_wire_3[493]),.i2(intermediate_wire_3[492]),.o(intermediate_reg_3[246])); 
xor_module xor_module_inst_3_578(.clk(clk),.reset(reset),.i1(intermediate_wire_3[491]),.i2(intermediate_wire_3[490]),.o(intermediate_reg_3[245])); 
xor_module xor_module_inst_3_579(.clk(clk),.reset(reset),.i1(intermediate_wire_3[489]),.i2(intermediate_wire_3[488]),.o(intermediate_reg_3[244])); 
xor_module xor_module_inst_3_580(.clk(clk),.reset(reset),.i1(intermediate_wire_3[487]),.i2(intermediate_wire_3[486]),.o(intermediate_reg_3[243])); 
xor_module xor_module_inst_3_581(.clk(clk),.reset(reset),.i1(intermediate_wire_3[485]),.i2(intermediate_wire_3[484]),.o(intermediate_reg_3[242])); 
mux_module mux_module_inst_3_582(.clk(clk),.reset(reset),.i1(intermediate_wire_3[483]),.i2(intermediate_wire_3[482]),.o(intermediate_reg_3[241]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_583(.clk(clk),.reset(reset),.i1(intermediate_wire_3[481]),.i2(intermediate_wire_3[480]),.o(intermediate_reg_3[240]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_584(.clk(clk),.reset(reset),.i1(intermediate_wire_3[479]),.i2(intermediate_wire_3[478]),.o(intermediate_reg_3[239]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_585(.clk(clk),.reset(reset),.i1(intermediate_wire_3[477]),.i2(intermediate_wire_3[476]),.o(intermediate_reg_3[238])); 
xor_module xor_module_inst_3_586(.clk(clk),.reset(reset),.i1(intermediate_wire_3[475]),.i2(intermediate_wire_3[474]),.o(intermediate_reg_3[237])); 
xor_module xor_module_inst_3_587(.clk(clk),.reset(reset),.i1(intermediate_wire_3[473]),.i2(intermediate_wire_3[472]),.o(intermediate_reg_3[236])); 
mux_module mux_module_inst_3_588(.clk(clk),.reset(reset),.i1(intermediate_wire_3[471]),.i2(intermediate_wire_3[470]),.o(intermediate_reg_3[235]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_589(.clk(clk),.reset(reset),.i1(intermediate_wire_3[469]),.i2(intermediate_wire_3[468]),.o(intermediate_reg_3[234]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_590(.clk(clk),.reset(reset),.i1(intermediate_wire_3[467]),.i2(intermediate_wire_3[466]),.o(intermediate_reg_3[233]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_591(.clk(clk),.reset(reset),.i1(intermediate_wire_3[465]),.i2(intermediate_wire_3[464]),.o(intermediate_reg_3[232])); 
mux_module mux_module_inst_3_592(.clk(clk),.reset(reset),.i1(intermediate_wire_3[463]),.i2(intermediate_wire_3[462]),.o(intermediate_reg_3[231]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_593(.clk(clk),.reset(reset),.i1(intermediate_wire_3[461]),.i2(intermediate_wire_3[460]),.o(intermediate_reg_3[230]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_594(.clk(clk),.reset(reset),.i1(intermediate_wire_3[459]),.i2(intermediate_wire_3[458]),.o(intermediate_reg_3[229])); 
xor_module xor_module_inst_3_595(.clk(clk),.reset(reset),.i1(intermediate_wire_3[457]),.i2(intermediate_wire_3[456]),.o(intermediate_reg_3[228])); 
mux_module mux_module_inst_3_596(.clk(clk),.reset(reset),.i1(intermediate_wire_3[455]),.i2(intermediate_wire_3[454]),.o(intermediate_reg_3[227]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_597(.clk(clk),.reset(reset),.i1(intermediate_wire_3[453]),.i2(intermediate_wire_3[452]),.o(intermediate_reg_3[226])); 
mux_module mux_module_inst_3_598(.clk(clk),.reset(reset),.i1(intermediate_wire_3[451]),.i2(intermediate_wire_3[450]),.o(intermediate_reg_3[225]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_599(.clk(clk),.reset(reset),.i1(intermediate_wire_3[449]),.i2(intermediate_wire_3[448]),.o(intermediate_reg_3[224]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_600(.clk(clk),.reset(reset),.i1(intermediate_wire_3[447]),.i2(intermediate_wire_3[446]),.o(intermediate_reg_3[223]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_601(.clk(clk),.reset(reset),.i1(intermediate_wire_3[445]),.i2(intermediate_wire_3[444]),.o(intermediate_reg_3[222]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_602(.clk(clk),.reset(reset),.i1(intermediate_wire_3[443]),.i2(intermediate_wire_3[442]),.o(intermediate_reg_3[221]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_603(.clk(clk),.reset(reset),.i1(intermediate_wire_3[441]),.i2(intermediate_wire_3[440]),.o(intermediate_reg_3[220]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_604(.clk(clk),.reset(reset),.i1(intermediate_wire_3[439]),.i2(intermediate_wire_3[438]),.o(intermediate_reg_3[219])); 
xor_module xor_module_inst_3_605(.clk(clk),.reset(reset),.i1(intermediate_wire_3[437]),.i2(intermediate_wire_3[436]),.o(intermediate_reg_3[218])); 
xor_module xor_module_inst_3_606(.clk(clk),.reset(reset),.i1(intermediate_wire_3[435]),.i2(intermediate_wire_3[434]),.o(intermediate_reg_3[217])); 
mux_module mux_module_inst_3_607(.clk(clk),.reset(reset),.i1(intermediate_wire_3[433]),.i2(intermediate_wire_3[432]),.o(intermediate_reg_3[216]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_608(.clk(clk),.reset(reset),.i1(intermediate_wire_3[431]),.i2(intermediate_wire_3[430]),.o(intermediate_reg_3[215])); 
xor_module xor_module_inst_3_609(.clk(clk),.reset(reset),.i1(intermediate_wire_3[429]),.i2(intermediate_wire_3[428]),.o(intermediate_reg_3[214])); 
mux_module mux_module_inst_3_610(.clk(clk),.reset(reset),.i1(intermediate_wire_3[427]),.i2(intermediate_wire_3[426]),.o(intermediate_reg_3[213]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_611(.clk(clk),.reset(reset),.i1(intermediate_wire_3[425]),.i2(intermediate_wire_3[424]),.o(intermediate_reg_3[212]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_612(.clk(clk),.reset(reset),.i1(intermediate_wire_3[423]),.i2(intermediate_wire_3[422]),.o(intermediate_reg_3[211])); 
mux_module mux_module_inst_3_613(.clk(clk),.reset(reset),.i1(intermediate_wire_3[421]),.i2(intermediate_wire_3[420]),.o(intermediate_reg_3[210]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_614(.clk(clk),.reset(reset),.i1(intermediate_wire_3[419]),.i2(intermediate_wire_3[418]),.o(intermediate_reg_3[209])); 
mux_module mux_module_inst_3_615(.clk(clk),.reset(reset),.i1(intermediate_wire_3[417]),.i2(intermediate_wire_3[416]),.o(intermediate_reg_3[208]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_616(.clk(clk),.reset(reset),.i1(intermediate_wire_3[415]),.i2(intermediate_wire_3[414]),.o(intermediate_reg_3[207])); 
mux_module mux_module_inst_3_617(.clk(clk),.reset(reset),.i1(intermediate_wire_3[413]),.i2(intermediate_wire_3[412]),.o(intermediate_reg_3[206]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_618(.clk(clk),.reset(reset),.i1(intermediate_wire_3[411]),.i2(intermediate_wire_3[410]),.o(intermediate_reg_3[205])); 
mux_module mux_module_inst_3_619(.clk(clk),.reset(reset),.i1(intermediate_wire_3[409]),.i2(intermediate_wire_3[408]),.o(intermediate_reg_3[204]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_620(.clk(clk),.reset(reset),.i1(intermediate_wire_3[407]),.i2(intermediate_wire_3[406]),.o(intermediate_reg_3[203]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_621(.clk(clk),.reset(reset),.i1(intermediate_wire_3[405]),.i2(intermediate_wire_3[404]),.o(intermediate_reg_3[202]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_622(.clk(clk),.reset(reset),.i1(intermediate_wire_3[403]),.i2(intermediate_wire_3[402]),.o(intermediate_reg_3[201]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_623(.clk(clk),.reset(reset),.i1(intermediate_wire_3[401]),.i2(intermediate_wire_3[400]),.o(intermediate_reg_3[200]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_624(.clk(clk),.reset(reset),.i1(intermediate_wire_3[399]),.i2(intermediate_wire_3[398]),.o(intermediate_reg_3[199]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_625(.clk(clk),.reset(reset),.i1(intermediate_wire_3[397]),.i2(intermediate_wire_3[396]),.o(intermediate_reg_3[198]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_626(.clk(clk),.reset(reset),.i1(intermediate_wire_3[395]),.i2(intermediate_wire_3[394]),.o(intermediate_reg_3[197])); 
mux_module mux_module_inst_3_627(.clk(clk),.reset(reset),.i1(intermediate_wire_3[393]),.i2(intermediate_wire_3[392]),.o(intermediate_reg_3[196]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_628(.clk(clk),.reset(reset),.i1(intermediate_wire_3[391]),.i2(intermediate_wire_3[390]),.o(intermediate_reg_3[195]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_629(.clk(clk),.reset(reset),.i1(intermediate_wire_3[389]),.i2(intermediate_wire_3[388]),.o(intermediate_reg_3[194])); 
xor_module xor_module_inst_3_630(.clk(clk),.reset(reset),.i1(intermediate_wire_3[387]),.i2(intermediate_wire_3[386]),.o(intermediate_reg_3[193])); 
xor_module xor_module_inst_3_631(.clk(clk),.reset(reset),.i1(intermediate_wire_3[385]),.i2(intermediate_wire_3[384]),.o(intermediate_reg_3[192])); 
mux_module mux_module_inst_3_632(.clk(clk),.reset(reset),.i1(intermediate_wire_3[383]),.i2(intermediate_wire_3[382]),.o(intermediate_reg_3[191]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_633(.clk(clk),.reset(reset),.i1(intermediate_wire_3[381]),.i2(intermediate_wire_3[380]),.o(intermediate_reg_3[190]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_634(.clk(clk),.reset(reset),.i1(intermediate_wire_3[379]),.i2(intermediate_wire_3[378]),.o(intermediate_reg_3[189])); 
xor_module xor_module_inst_3_635(.clk(clk),.reset(reset),.i1(intermediate_wire_3[377]),.i2(intermediate_wire_3[376]),.o(intermediate_reg_3[188])); 
xor_module xor_module_inst_3_636(.clk(clk),.reset(reset),.i1(intermediate_wire_3[375]),.i2(intermediate_wire_3[374]),.o(intermediate_reg_3[187])); 
xor_module xor_module_inst_3_637(.clk(clk),.reset(reset),.i1(intermediate_wire_3[373]),.i2(intermediate_wire_3[372]),.o(intermediate_reg_3[186])); 
mux_module mux_module_inst_3_638(.clk(clk),.reset(reset),.i1(intermediate_wire_3[371]),.i2(intermediate_wire_3[370]),.o(intermediate_reg_3[185]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_639(.clk(clk),.reset(reset),.i1(intermediate_wire_3[369]),.i2(intermediate_wire_3[368]),.o(intermediate_reg_3[184]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_640(.clk(clk),.reset(reset),.i1(intermediate_wire_3[367]),.i2(intermediate_wire_3[366]),.o(intermediate_reg_3[183])); 
xor_module xor_module_inst_3_641(.clk(clk),.reset(reset),.i1(intermediate_wire_3[365]),.i2(intermediate_wire_3[364]),.o(intermediate_reg_3[182])); 
xor_module xor_module_inst_3_642(.clk(clk),.reset(reset),.i1(intermediate_wire_3[363]),.i2(intermediate_wire_3[362]),.o(intermediate_reg_3[181])); 
xor_module xor_module_inst_3_643(.clk(clk),.reset(reset),.i1(intermediate_wire_3[361]),.i2(intermediate_wire_3[360]),.o(intermediate_reg_3[180])); 
mux_module mux_module_inst_3_644(.clk(clk),.reset(reset),.i1(intermediate_wire_3[359]),.i2(intermediate_wire_3[358]),.o(intermediate_reg_3[179]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_645(.clk(clk),.reset(reset),.i1(intermediate_wire_3[357]),.i2(intermediate_wire_3[356]),.o(intermediate_reg_3[178]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_646(.clk(clk),.reset(reset),.i1(intermediate_wire_3[355]),.i2(intermediate_wire_3[354]),.o(intermediate_reg_3[177])); 
mux_module mux_module_inst_3_647(.clk(clk),.reset(reset),.i1(intermediate_wire_3[353]),.i2(intermediate_wire_3[352]),.o(intermediate_reg_3[176]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_648(.clk(clk),.reset(reset),.i1(intermediate_wire_3[351]),.i2(intermediate_wire_3[350]),.o(intermediate_reg_3[175])); 
xor_module xor_module_inst_3_649(.clk(clk),.reset(reset),.i1(intermediate_wire_3[349]),.i2(intermediate_wire_3[348]),.o(intermediate_reg_3[174])); 
mux_module mux_module_inst_3_650(.clk(clk),.reset(reset),.i1(intermediate_wire_3[347]),.i2(intermediate_wire_3[346]),.o(intermediate_reg_3[173]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_651(.clk(clk),.reset(reset),.i1(intermediate_wire_3[345]),.i2(intermediate_wire_3[344]),.o(intermediate_reg_3[172])); 
mux_module mux_module_inst_3_652(.clk(clk),.reset(reset),.i1(intermediate_wire_3[343]),.i2(intermediate_wire_3[342]),.o(intermediate_reg_3[171]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_653(.clk(clk),.reset(reset),.i1(intermediate_wire_3[341]),.i2(intermediate_wire_3[340]),.o(intermediate_reg_3[170])); 
mux_module mux_module_inst_3_654(.clk(clk),.reset(reset),.i1(intermediate_wire_3[339]),.i2(intermediate_wire_3[338]),.o(intermediate_reg_3[169]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_655(.clk(clk),.reset(reset),.i1(intermediate_wire_3[337]),.i2(intermediate_wire_3[336]),.o(intermediate_reg_3[168]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_656(.clk(clk),.reset(reset),.i1(intermediate_wire_3[335]),.i2(intermediate_wire_3[334]),.o(intermediate_reg_3[167]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_657(.clk(clk),.reset(reset),.i1(intermediate_wire_3[333]),.i2(intermediate_wire_3[332]),.o(intermediate_reg_3[166]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_658(.clk(clk),.reset(reset),.i1(intermediate_wire_3[331]),.i2(intermediate_wire_3[330]),.o(intermediate_reg_3[165]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_659(.clk(clk),.reset(reset),.i1(intermediate_wire_3[329]),.i2(intermediate_wire_3[328]),.o(intermediate_reg_3[164]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_660(.clk(clk),.reset(reset),.i1(intermediate_wire_3[327]),.i2(intermediate_wire_3[326]),.o(intermediate_reg_3[163])); 
xor_module xor_module_inst_3_661(.clk(clk),.reset(reset),.i1(intermediate_wire_3[325]),.i2(intermediate_wire_3[324]),.o(intermediate_reg_3[162])); 
mux_module mux_module_inst_3_662(.clk(clk),.reset(reset),.i1(intermediate_wire_3[323]),.i2(intermediate_wire_3[322]),.o(intermediate_reg_3[161]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_663(.clk(clk),.reset(reset),.i1(intermediate_wire_3[321]),.i2(intermediate_wire_3[320]),.o(intermediate_reg_3[160])); 
xor_module xor_module_inst_3_664(.clk(clk),.reset(reset),.i1(intermediate_wire_3[319]),.i2(intermediate_wire_3[318]),.o(intermediate_reg_3[159])); 
mux_module mux_module_inst_3_665(.clk(clk),.reset(reset),.i1(intermediate_wire_3[317]),.i2(intermediate_wire_3[316]),.o(intermediate_reg_3[158]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_666(.clk(clk),.reset(reset),.i1(intermediate_wire_3[315]),.i2(intermediate_wire_3[314]),.o(intermediate_reg_3[157])); 
mux_module mux_module_inst_3_667(.clk(clk),.reset(reset),.i1(intermediate_wire_3[313]),.i2(intermediate_wire_3[312]),.o(intermediate_reg_3[156]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_668(.clk(clk),.reset(reset),.i1(intermediate_wire_3[311]),.i2(intermediate_wire_3[310]),.o(intermediate_reg_3[155])); 
mux_module mux_module_inst_3_669(.clk(clk),.reset(reset),.i1(intermediate_wire_3[309]),.i2(intermediate_wire_3[308]),.o(intermediate_reg_3[154]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_670(.clk(clk),.reset(reset),.i1(intermediate_wire_3[307]),.i2(intermediate_wire_3[306]),.o(intermediate_reg_3[153])); 
mux_module mux_module_inst_3_671(.clk(clk),.reset(reset),.i1(intermediate_wire_3[305]),.i2(intermediate_wire_3[304]),.o(intermediate_reg_3[152]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_672(.clk(clk),.reset(reset),.i1(intermediate_wire_3[303]),.i2(intermediate_wire_3[302]),.o(intermediate_reg_3[151]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_673(.clk(clk),.reset(reset),.i1(intermediate_wire_3[301]),.i2(intermediate_wire_3[300]),.o(intermediate_reg_3[150]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_674(.clk(clk),.reset(reset),.i1(intermediate_wire_3[299]),.i2(intermediate_wire_3[298]),.o(intermediate_reg_3[149]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_675(.clk(clk),.reset(reset),.i1(intermediate_wire_3[297]),.i2(intermediate_wire_3[296]),.o(intermediate_reg_3[148])); 
xor_module xor_module_inst_3_676(.clk(clk),.reset(reset),.i1(intermediate_wire_3[295]),.i2(intermediate_wire_3[294]),.o(intermediate_reg_3[147])); 
mux_module mux_module_inst_3_677(.clk(clk),.reset(reset),.i1(intermediate_wire_3[293]),.i2(intermediate_wire_3[292]),.o(intermediate_reg_3[146]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_678(.clk(clk),.reset(reset),.i1(intermediate_wire_3[291]),.i2(intermediate_wire_3[290]),.o(intermediate_reg_3[145])); 
mux_module mux_module_inst_3_679(.clk(clk),.reset(reset),.i1(intermediate_wire_3[289]),.i2(intermediate_wire_3[288]),.o(intermediate_reg_3[144]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_680(.clk(clk),.reset(reset),.i1(intermediate_wire_3[287]),.i2(intermediate_wire_3[286]),.o(intermediate_reg_3[143])); 
mux_module mux_module_inst_3_681(.clk(clk),.reset(reset),.i1(intermediate_wire_3[285]),.i2(intermediate_wire_3[284]),.o(intermediate_reg_3[142]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_682(.clk(clk),.reset(reset),.i1(intermediate_wire_3[283]),.i2(intermediate_wire_3[282]),.o(intermediate_reg_3[141]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_683(.clk(clk),.reset(reset),.i1(intermediate_wire_3[281]),.i2(intermediate_wire_3[280]),.o(intermediate_reg_3[140])); 
mux_module mux_module_inst_3_684(.clk(clk),.reset(reset),.i1(intermediate_wire_3[279]),.i2(intermediate_wire_3[278]),.o(intermediate_reg_3[139]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_685(.clk(clk),.reset(reset),.i1(intermediate_wire_3[277]),.i2(intermediate_wire_3[276]),.o(intermediate_reg_3[138])); 
mux_module mux_module_inst_3_686(.clk(clk),.reset(reset),.i1(intermediate_wire_3[275]),.i2(intermediate_wire_3[274]),.o(intermediate_reg_3[137]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_687(.clk(clk),.reset(reset),.i1(intermediate_wire_3[273]),.i2(intermediate_wire_3[272]),.o(intermediate_reg_3[136])); 
mux_module mux_module_inst_3_688(.clk(clk),.reset(reset),.i1(intermediate_wire_3[271]),.i2(intermediate_wire_3[270]),.o(intermediate_reg_3[135]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_689(.clk(clk),.reset(reset),.i1(intermediate_wire_3[269]),.i2(intermediate_wire_3[268]),.o(intermediate_reg_3[134])); 
mux_module mux_module_inst_3_690(.clk(clk),.reset(reset),.i1(intermediate_wire_3[267]),.i2(intermediate_wire_3[266]),.o(intermediate_reg_3[133]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_691(.clk(clk),.reset(reset),.i1(intermediate_wire_3[265]),.i2(intermediate_wire_3[264]),.o(intermediate_reg_3[132]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_692(.clk(clk),.reset(reset),.i1(intermediate_wire_3[263]),.i2(intermediate_wire_3[262]),.o(intermediate_reg_3[131])); 
xor_module xor_module_inst_3_693(.clk(clk),.reset(reset),.i1(intermediate_wire_3[261]),.i2(intermediate_wire_3[260]),.o(intermediate_reg_3[130])); 
xor_module xor_module_inst_3_694(.clk(clk),.reset(reset),.i1(intermediate_wire_3[259]),.i2(intermediate_wire_3[258]),.o(intermediate_reg_3[129])); 
xor_module xor_module_inst_3_695(.clk(clk),.reset(reset),.i1(intermediate_wire_3[257]),.i2(intermediate_wire_3[256]),.o(intermediate_reg_3[128])); 
xor_module xor_module_inst_3_696(.clk(clk),.reset(reset),.i1(intermediate_wire_3[255]),.i2(intermediate_wire_3[254]),.o(intermediate_reg_3[127])); 
xor_module xor_module_inst_3_697(.clk(clk),.reset(reset),.i1(intermediate_wire_3[253]),.i2(intermediate_wire_3[252]),.o(intermediate_reg_3[126])); 
mux_module mux_module_inst_3_698(.clk(clk),.reset(reset),.i1(intermediate_wire_3[251]),.i2(intermediate_wire_3[250]),.o(intermediate_reg_3[125]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_699(.clk(clk),.reset(reset),.i1(intermediate_wire_3[249]),.i2(intermediate_wire_3[248]),.o(intermediate_reg_3[124]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_700(.clk(clk),.reset(reset),.i1(intermediate_wire_3[247]),.i2(intermediate_wire_3[246]),.o(intermediate_reg_3[123]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_701(.clk(clk),.reset(reset),.i1(intermediate_wire_3[245]),.i2(intermediate_wire_3[244]),.o(intermediate_reg_3[122]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_702(.clk(clk),.reset(reset),.i1(intermediate_wire_3[243]),.i2(intermediate_wire_3[242]),.o(intermediate_reg_3[121])); 
mux_module mux_module_inst_3_703(.clk(clk),.reset(reset),.i1(intermediate_wire_3[241]),.i2(intermediate_wire_3[240]),.o(intermediate_reg_3[120]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_704(.clk(clk),.reset(reset),.i1(intermediate_wire_3[239]),.i2(intermediate_wire_3[238]),.o(intermediate_reg_3[119])); 
mux_module mux_module_inst_3_705(.clk(clk),.reset(reset),.i1(intermediate_wire_3[237]),.i2(intermediate_wire_3[236]),.o(intermediate_reg_3[118]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_706(.clk(clk),.reset(reset),.i1(intermediate_wire_3[235]),.i2(intermediate_wire_3[234]),.o(intermediate_reg_3[117])); 
mux_module mux_module_inst_3_707(.clk(clk),.reset(reset),.i1(intermediate_wire_3[233]),.i2(intermediate_wire_3[232]),.o(intermediate_reg_3[116]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_708(.clk(clk),.reset(reset),.i1(intermediate_wire_3[231]),.i2(intermediate_wire_3[230]),.o(intermediate_reg_3[115])); 
mux_module mux_module_inst_3_709(.clk(clk),.reset(reset),.i1(intermediate_wire_3[229]),.i2(intermediate_wire_3[228]),.o(intermediate_reg_3[114]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_710(.clk(clk),.reset(reset),.i1(intermediate_wire_3[227]),.i2(intermediate_wire_3[226]),.o(intermediate_reg_3[113])); 
mux_module mux_module_inst_3_711(.clk(clk),.reset(reset),.i1(intermediate_wire_3[225]),.i2(intermediate_wire_3[224]),.o(intermediate_reg_3[112]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_712(.clk(clk),.reset(reset),.i1(intermediate_wire_3[223]),.i2(intermediate_wire_3[222]),.o(intermediate_reg_3[111]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_713(.clk(clk),.reset(reset),.i1(intermediate_wire_3[221]),.i2(intermediate_wire_3[220]),.o(intermediate_reg_3[110])); 
mux_module mux_module_inst_3_714(.clk(clk),.reset(reset),.i1(intermediate_wire_3[219]),.i2(intermediate_wire_3[218]),.o(intermediate_reg_3[109]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_715(.clk(clk),.reset(reset),.i1(intermediate_wire_3[217]),.i2(intermediate_wire_3[216]),.o(intermediate_reg_3[108])); 
mux_module mux_module_inst_3_716(.clk(clk),.reset(reset),.i1(intermediate_wire_3[215]),.i2(intermediate_wire_3[214]),.o(intermediate_reg_3[107]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_717(.clk(clk),.reset(reset),.i1(intermediate_wire_3[213]),.i2(intermediate_wire_3[212]),.o(intermediate_reg_3[106])); 
mux_module mux_module_inst_3_718(.clk(clk),.reset(reset),.i1(intermediate_wire_3[211]),.i2(intermediate_wire_3[210]),.o(intermediate_reg_3[105]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_719(.clk(clk),.reset(reset),.i1(intermediate_wire_3[209]),.i2(intermediate_wire_3[208]),.o(intermediate_reg_3[104])); 
mux_module mux_module_inst_3_720(.clk(clk),.reset(reset),.i1(intermediate_wire_3[207]),.i2(intermediate_wire_3[206]),.o(intermediate_reg_3[103]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_721(.clk(clk),.reset(reset),.i1(intermediate_wire_3[205]),.i2(intermediate_wire_3[204]),.o(intermediate_reg_3[102])); 
xor_module xor_module_inst_3_722(.clk(clk),.reset(reset),.i1(intermediate_wire_3[203]),.i2(intermediate_wire_3[202]),.o(intermediate_reg_3[101])); 
mux_module mux_module_inst_3_723(.clk(clk),.reset(reset),.i1(intermediate_wire_3[201]),.i2(intermediate_wire_3[200]),.o(intermediate_reg_3[100]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_724(.clk(clk),.reset(reset),.i1(intermediate_wire_3[199]),.i2(intermediate_wire_3[198]),.o(intermediate_reg_3[99]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_725(.clk(clk),.reset(reset),.i1(intermediate_wire_3[197]),.i2(intermediate_wire_3[196]),.o(intermediate_reg_3[98]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_726(.clk(clk),.reset(reset),.i1(intermediate_wire_3[195]),.i2(intermediate_wire_3[194]),.o(intermediate_reg_3[97])); 
xor_module xor_module_inst_3_727(.clk(clk),.reset(reset),.i1(intermediate_wire_3[193]),.i2(intermediate_wire_3[192]),.o(intermediate_reg_3[96])); 
xor_module xor_module_inst_3_728(.clk(clk),.reset(reset),.i1(intermediate_wire_3[191]),.i2(intermediate_wire_3[190]),.o(intermediate_reg_3[95])); 
mux_module mux_module_inst_3_729(.clk(clk),.reset(reset),.i1(intermediate_wire_3[189]),.i2(intermediate_wire_3[188]),.o(intermediate_reg_3[94]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_730(.clk(clk),.reset(reset),.i1(intermediate_wire_3[187]),.i2(intermediate_wire_3[186]),.o(intermediate_reg_3[93]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_731(.clk(clk),.reset(reset),.i1(intermediate_wire_3[185]),.i2(intermediate_wire_3[184]),.o(intermediate_reg_3[92])); 
xor_module xor_module_inst_3_732(.clk(clk),.reset(reset),.i1(intermediate_wire_3[183]),.i2(intermediate_wire_3[182]),.o(intermediate_reg_3[91])); 
mux_module mux_module_inst_3_733(.clk(clk),.reset(reset),.i1(intermediate_wire_3[181]),.i2(intermediate_wire_3[180]),.o(intermediate_reg_3[90]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_734(.clk(clk),.reset(reset),.i1(intermediate_wire_3[179]),.i2(intermediate_wire_3[178]),.o(intermediate_reg_3[89]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_735(.clk(clk),.reset(reset),.i1(intermediate_wire_3[177]),.i2(intermediate_wire_3[176]),.o(intermediate_reg_3[88]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_736(.clk(clk),.reset(reset),.i1(intermediate_wire_3[175]),.i2(intermediate_wire_3[174]),.o(intermediate_reg_3[87])); 
xor_module xor_module_inst_3_737(.clk(clk),.reset(reset),.i1(intermediate_wire_3[173]),.i2(intermediate_wire_3[172]),.o(intermediate_reg_3[86])); 
xor_module xor_module_inst_3_738(.clk(clk),.reset(reset),.i1(intermediate_wire_3[171]),.i2(intermediate_wire_3[170]),.o(intermediate_reg_3[85])); 
xor_module xor_module_inst_3_739(.clk(clk),.reset(reset),.i1(intermediate_wire_3[169]),.i2(intermediate_wire_3[168]),.o(intermediate_reg_3[84])); 
mux_module mux_module_inst_3_740(.clk(clk),.reset(reset),.i1(intermediate_wire_3[167]),.i2(intermediate_wire_3[166]),.o(intermediate_reg_3[83]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_741(.clk(clk),.reset(reset),.i1(intermediate_wire_3[165]),.i2(intermediate_wire_3[164]),.o(intermediate_reg_3[82]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_742(.clk(clk),.reset(reset),.i1(intermediate_wire_3[163]),.i2(intermediate_wire_3[162]),.o(intermediate_reg_3[81]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_743(.clk(clk),.reset(reset),.i1(intermediate_wire_3[161]),.i2(intermediate_wire_3[160]),.o(intermediate_reg_3[80])); 
xor_module xor_module_inst_3_744(.clk(clk),.reset(reset),.i1(intermediate_wire_3[159]),.i2(intermediate_wire_3[158]),.o(intermediate_reg_3[79])); 
mux_module mux_module_inst_3_745(.clk(clk),.reset(reset),.i1(intermediate_wire_3[157]),.i2(intermediate_wire_3[156]),.o(intermediate_reg_3[78]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_746(.clk(clk),.reset(reset),.i1(intermediate_wire_3[155]),.i2(intermediate_wire_3[154]),.o(intermediate_reg_3[77]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_747(.clk(clk),.reset(reset),.i1(intermediate_wire_3[153]),.i2(intermediate_wire_3[152]),.o(intermediate_reg_3[76]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_748(.clk(clk),.reset(reset),.i1(intermediate_wire_3[151]),.i2(intermediate_wire_3[150]),.o(intermediate_reg_3[75])); 
mux_module mux_module_inst_3_749(.clk(clk),.reset(reset),.i1(intermediate_wire_3[149]),.i2(intermediate_wire_3[148]),.o(intermediate_reg_3[74]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_750(.clk(clk),.reset(reset),.i1(intermediate_wire_3[147]),.i2(intermediate_wire_3[146]),.o(intermediate_reg_3[73])); 
xor_module xor_module_inst_3_751(.clk(clk),.reset(reset),.i1(intermediate_wire_3[145]),.i2(intermediate_wire_3[144]),.o(intermediate_reg_3[72])); 
mux_module mux_module_inst_3_752(.clk(clk),.reset(reset),.i1(intermediate_wire_3[143]),.i2(intermediate_wire_3[142]),.o(intermediate_reg_3[71]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_753(.clk(clk),.reset(reset),.i1(intermediate_wire_3[141]),.i2(intermediate_wire_3[140]),.o(intermediate_reg_3[70]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_754(.clk(clk),.reset(reset),.i1(intermediate_wire_3[139]),.i2(intermediate_wire_3[138]),.o(intermediate_reg_3[69])); 
mux_module mux_module_inst_3_755(.clk(clk),.reset(reset),.i1(intermediate_wire_3[137]),.i2(intermediate_wire_3[136]),.o(intermediate_reg_3[68]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_756(.clk(clk),.reset(reset),.i1(intermediate_wire_3[135]),.i2(intermediate_wire_3[134]),.o(intermediate_reg_3[67])); 
xor_module xor_module_inst_3_757(.clk(clk),.reset(reset),.i1(intermediate_wire_3[133]),.i2(intermediate_wire_3[132]),.o(intermediate_reg_3[66])); 
xor_module xor_module_inst_3_758(.clk(clk),.reset(reset),.i1(intermediate_wire_3[131]),.i2(intermediate_wire_3[130]),.o(intermediate_reg_3[65])); 
mux_module mux_module_inst_3_759(.clk(clk),.reset(reset),.i1(intermediate_wire_3[129]),.i2(intermediate_wire_3[128]),.o(intermediate_reg_3[64]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_760(.clk(clk),.reset(reset),.i1(intermediate_wire_3[127]),.i2(intermediate_wire_3[126]),.o(intermediate_reg_3[63]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_761(.clk(clk),.reset(reset),.i1(intermediate_wire_3[125]),.i2(intermediate_wire_3[124]),.o(intermediate_reg_3[62]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_762(.clk(clk),.reset(reset),.i1(intermediate_wire_3[123]),.i2(intermediate_wire_3[122]),.o(intermediate_reg_3[61]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_763(.clk(clk),.reset(reset),.i1(intermediate_wire_3[121]),.i2(intermediate_wire_3[120]),.o(intermediate_reg_3[60]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_764(.clk(clk),.reset(reset),.i1(intermediate_wire_3[119]),.i2(intermediate_wire_3[118]),.o(intermediate_reg_3[59]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_765(.clk(clk),.reset(reset),.i1(intermediate_wire_3[117]),.i2(intermediate_wire_3[116]),.o(intermediate_reg_3[58])); 
mux_module mux_module_inst_3_766(.clk(clk),.reset(reset),.i1(intermediate_wire_3[115]),.i2(intermediate_wire_3[114]),.o(intermediate_reg_3[57]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_767(.clk(clk),.reset(reset),.i1(intermediate_wire_3[113]),.i2(intermediate_wire_3[112]),.o(intermediate_reg_3[56])); 
mux_module mux_module_inst_3_768(.clk(clk),.reset(reset),.i1(intermediate_wire_3[111]),.i2(intermediate_wire_3[110]),.o(intermediate_reg_3[55]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_769(.clk(clk),.reset(reset),.i1(intermediate_wire_3[109]),.i2(intermediate_wire_3[108]),.o(intermediate_reg_3[54]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_770(.clk(clk),.reset(reset),.i1(intermediate_wire_3[107]),.i2(intermediate_wire_3[106]),.o(intermediate_reg_3[53])); 
mux_module mux_module_inst_3_771(.clk(clk),.reset(reset),.i1(intermediate_wire_3[105]),.i2(intermediate_wire_3[104]),.o(intermediate_reg_3[52]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_772(.clk(clk),.reset(reset),.i1(intermediate_wire_3[103]),.i2(intermediate_wire_3[102]),.o(intermediate_reg_3[51])); 
xor_module xor_module_inst_3_773(.clk(clk),.reset(reset),.i1(intermediate_wire_3[101]),.i2(intermediate_wire_3[100]),.o(intermediate_reg_3[50])); 
xor_module xor_module_inst_3_774(.clk(clk),.reset(reset),.i1(intermediate_wire_3[99]),.i2(intermediate_wire_3[98]),.o(intermediate_reg_3[49])); 
mux_module mux_module_inst_3_775(.clk(clk),.reset(reset),.i1(intermediate_wire_3[97]),.i2(intermediate_wire_3[96]),.o(intermediate_reg_3[48]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_776(.clk(clk),.reset(reset),.i1(intermediate_wire_3[95]),.i2(intermediate_wire_3[94]),.o(intermediate_reg_3[47]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_777(.clk(clk),.reset(reset),.i1(intermediate_wire_3[93]),.i2(intermediate_wire_3[92]),.o(intermediate_reg_3[46])); 
xor_module xor_module_inst_3_778(.clk(clk),.reset(reset),.i1(intermediate_wire_3[91]),.i2(intermediate_wire_3[90]),.o(intermediate_reg_3[45])); 
xor_module xor_module_inst_3_779(.clk(clk),.reset(reset),.i1(intermediate_wire_3[89]),.i2(intermediate_wire_3[88]),.o(intermediate_reg_3[44])); 
mux_module mux_module_inst_3_780(.clk(clk),.reset(reset),.i1(intermediate_wire_3[87]),.i2(intermediate_wire_3[86]),.o(intermediate_reg_3[43]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_781(.clk(clk),.reset(reset),.i1(intermediate_wire_3[85]),.i2(intermediate_wire_3[84]),.o(intermediate_reg_3[42]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_782(.clk(clk),.reset(reset),.i1(intermediate_wire_3[83]),.i2(intermediate_wire_3[82]),.o(intermediate_reg_3[41]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_783(.clk(clk),.reset(reset),.i1(intermediate_wire_3[81]),.i2(intermediate_wire_3[80]),.o(intermediate_reg_3[40]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_784(.clk(clk),.reset(reset),.i1(intermediate_wire_3[79]),.i2(intermediate_wire_3[78]),.o(intermediate_reg_3[39]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_785(.clk(clk),.reset(reset),.i1(intermediate_wire_3[77]),.i2(intermediate_wire_3[76]),.o(intermediate_reg_3[38]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_786(.clk(clk),.reset(reset),.i1(intermediate_wire_3[75]),.i2(intermediate_wire_3[74]),.o(intermediate_reg_3[37])); 
mux_module mux_module_inst_3_787(.clk(clk),.reset(reset),.i1(intermediate_wire_3[73]),.i2(intermediate_wire_3[72]),.o(intermediate_reg_3[36]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_788(.clk(clk),.reset(reset),.i1(intermediate_wire_3[71]),.i2(intermediate_wire_3[70]),.o(intermediate_reg_3[35]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_789(.clk(clk),.reset(reset),.i1(intermediate_wire_3[69]),.i2(intermediate_wire_3[68]),.o(intermediate_reg_3[34])); 
xor_module xor_module_inst_3_790(.clk(clk),.reset(reset),.i1(intermediate_wire_3[67]),.i2(intermediate_wire_3[66]),.o(intermediate_reg_3[33])); 
mux_module mux_module_inst_3_791(.clk(clk),.reset(reset),.i1(intermediate_wire_3[65]),.i2(intermediate_wire_3[64]),.o(intermediate_reg_3[32]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_792(.clk(clk),.reset(reset),.i1(intermediate_wire_3[63]),.i2(intermediate_wire_3[62]),.o(intermediate_reg_3[31]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_793(.clk(clk),.reset(reset),.i1(intermediate_wire_3[61]),.i2(intermediate_wire_3[60]),.o(intermediate_reg_3[30])); 
mux_module mux_module_inst_3_794(.clk(clk),.reset(reset),.i1(intermediate_wire_3[59]),.i2(intermediate_wire_3[58]),.o(intermediate_reg_3[29]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_795(.clk(clk),.reset(reset),.i1(intermediate_wire_3[57]),.i2(intermediate_wire_3[56]),.o(intermediate_reg_3[28])); 
mux_module mux_module_inst_3_796(.clk(clk),.reset(reset),.i1(intermediate_wire_3[55]),.i2(intermediate_wire_3[54]),.o(intermediate_reg_3[27]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_797(.clk(clk),.reset(reset),.i1(intermediate_wire_3[53]),.i2(intermediate_wire_3[52]),.o(intermediate_reg_3[26])); 
xor_module xor_module_inst_3_798(.clk(clk),.reset(reset),.i1(intermediate_wire_3[51]),.i2(intermediate_wire_3[50]),.o(intermediate_reg_3[25])); 
mux_module mux_module_inst_3_799(.clk(clk),.reset(reset),.i1(intermediate_wire_3[49]),.i2(intermediate_wire_3[48]),.o(intermediate_reg_3[24]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_800(.clk(clk),.reset(reset),.i1(intermediate_wire_3[47]),.i2(intermediate_wire_3[46]),.o(intermediate_reg_3[23])); 
mux_module mux_module_inst_3_801(.clk(clk),.reset(reset),.i1(intermediate_wire_3[45]),.i2(intermediate_wire_3[44]),.o(intermediate_reg_3[22]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_802(.clk(clk),.reset(reset),.i1(intermediate_wire_3[43]),.i2(intermediate_wire_3[42]),.o(intermediate_reg_3[21]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_803(.clk(clk),.reset(reset),.i1(intermediate_wire_3[41]),.i2(intermediate_wire_3[40]),.o(intermediate_reg_3[20]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_804(.clk(clk),.reset(reset),.i1(intermediate_wire_3[39]),.i2(intermediate_wire_3[38]),.o(intermediate_reg_3[19])); 
mux_module mux_module_inst_3_805(.clk(clk),.reset(reset),.i1(intermediate_wire_3[37]),.i2(intermediate_wire_3[36]),.o(intermediate_reg_3[18]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_806(.clk(clk),.reset(reset),.i1(intermediate_wire_3[35]),.i2(intermediate_wire_3[34]),.o(intermediate_reg_3[17])); 
xor_module xor_module_inst_3_807(.clk(clk),.reset(reset),.i1(intermediate_wire_3[33]),.i2(intermediate_wire_3[32]),.o(intermediate_reg_3[16])); 
mux_module mux_module_inst_3_808(.clk(clk),.reset(reset),.i1(intermediate_wire_3[31]),.i2(intermediate_wire_3[30]),.o(intermediate_reg_3[15]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_809(.clk(clk),.reset(reset),.i1(intermediate_wire_3[29]),.i2(intermediate_wire_3[28]),.o(intermediate_reg_3[14]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_810(.clk(clk),.reset(reset),.i1(intermediate_wire_3[27]),.i2(intermediate_wire_3[26]),.o(intermediate_reg_3[13])); 
xor_module xor_module_inst_3_811(.clk(clk),.reset(reset),.i1(intermediate_wire_3[25]),.i2(intermediate_wire_3[24]),.o(intermediate_reg_3[12])); 
mux_module mux_module_inst_3_812(.clk(clk),.reset(reset),.i1(intermediate_wire_3[23]),.i2(intermediate_wire_3[22]),.o(intermediate_reg_3[11]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_813(.clk(clk),.reset(reset),.i1(intermediate_wire_3[21]),.i2(intermediate_wire_3[20]),.o(intermediate_reg_3[10])); 
mux_module mux_module_inst_3_814(.clk(clk),.reset(reset),.i1(intermediate_wire_3[19]),.i2(intermediate_wire_3[18]),.o(intermediate_reg_3[9]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_815(.clk(clk),.reset(reset),.i1(intermediate_wire_3[17]),.i2(intermediate_wire_3[16]),.o(intermediate_reg_3[8]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_816(.clk(clk),.reset(reset),.i1(intermediate_wire_3[15]),.i2(intermediate_wire_3[14]),.o(intermediate_reg_3[7])); 
xor_module xor_module_inst_3_817(.clk(clk),.reset(reset),.i1(intermediate_wire_3[13]),.i2(intermediate_wire_3[12]),.o(intermediate_reg_3[6])); 
mux_module mux_module_inst_3_818(.clk(clk),.reset(reset),.i1(intermediate_wire_3[11]),.i2(intermediate_wire_3[10]),.o(intermediate_reg_3[5]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_819(.clk(clk),.reset(reset),.i1(intermediate_wire_3[9]),.i2(intermediate_wire_3[8]),.o(intermediate_reg_3[4]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_820(.clk(clk),.reset(reset),.i1(intermediate_wire_3[7]),.i2(intermediate_wire_3[6]),.o(intermediate_reg_3[3]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_821(.clk(clk),.reset(reset),.i1(intermediate_wire_3[5]),.i2(intermediate_wire_3[4]),.o(intermediate_reg_3[2]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_822(.clk(clk),.reset(reset),.i1(intermediate_wire_3[3]),.i2(intermediate_wire_3[2]),.o(intermediate_reg_3[1]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_823(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1]),.i2(intermediate_wire_3[0]),.o(intermediate_reg_3[0]),.sel(intermediate_reg_2[0])); 
always@(posedge clk) begin 
outp [823:0] <= intermediate_reg_3; 
outp[835:824] <= intermediate_reg_3[11:0] ; 
end 
endmodule 
 

module interface_14(input [119:0] inp, output reg [417:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[119:0] <= inp ; 
outp[239:120] <= inp ; 
outp[359:240] <= inp ; 
outp[417:360] <= inp[57:0] ; 
end 
endmodule 

module interface_15(input [223:0] inp, output reg [127:0] outp, input clk, input reset);
reg [223:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
wire [111:0]intermediate_reg_1; 
 
xor_module xor_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
xor_module xor_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
xor_module xor_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
mux_module mux_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
mux_module mux_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
xor_module xor_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
xor_module xor_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
xor_module xor_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
xor_module xor_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
xor_module xor_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
xor_module xor_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
xor_module xor_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
mux_module mux_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
xor_module xor_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
xor_module xor_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
mux_module mux_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
mux_module mux_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
xor_module xor_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [111:0] <= intermediate_reg_1; 
outp[127:112] <= intermediate_reg_1[15:0] ; 
end 
endmodule 
 

module interface_16(input [119:0] inp, output reg [383:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[119:0] <= inp ; 
outp[239:120] <= inp ; 
outp[359:240] <= inp ; 
outp[383:360] <= inp[23:0] ; 
end 
endmodule 

module interface_17(input [863:0] inp, output reg [1151:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[863:0] <= inp ; 
outp[1151:864] <= inp[287:0] ; 
end 
endmodule 

module dbram_2048_40bit_module_2(input clk, input reset, input[207:0] inp, output [159:0] outp); 

dbram_2048_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[103:0]),.outp(outp[79:0])); 

dbram_2048_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[207:104]),.outp(outp[159:80])); 

endmodule 

module systolic_array_4_fp16bit_2(input clk, input reset, input[835:0] inp, output [447:0] outp); 

systolic_array_4_fp16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[417:0]),.outp(outp[223:0])); 

systolic_array_4_fp16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[835:418]),.outp(outp[447:224])); 

endmodule 

module dbram_2048_60bit_module_12(input clk, input reset, input[1727:0] inp, output [1439:0] outp); 

dbram_2048_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[143:0]),.outp(outp[119:0])); 

dbram_2048_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[287:144]),.outp(outp[239:120])); 

dbram_2048_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[431:288]),.outp(outp[359:240])); 

dbram_2048_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[575:432]),.outp(outp[479:360])); 

dbram_2048_60bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[719:576]),.outp(outp[599:480])); 

dbram_2048_60bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[863:720]),.outp(outp[719:600])); 

dbram_2048_60bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1007:864]),.outp(outp[839:720])); 

dbram_2048_60bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[1151:1008]),.outp(outp[959:840])); 

dbram_2048_60bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[1295:1152]),.outp(outp[1079:960])); 

dbram_2048_60bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1439:1296]),.outp(outp[1199:1080])); 

dbram_2048_60bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[1583:1440]),.outp(outp[1319:1200])); 

dbram_2048_60bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[1727:1584]),.outp(outp[1439:1320])); 

endmodule 

module dbram_4096_40bit_module_10(input clk, input reset, input[1059:0] inp, output [799:0] outp); 

dbram_4096_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[105:0]),.outp(outp[79:0])); 

dbram_4096_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[211:106]),.outp(outp[159:80])); 

dbram_4096_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[317:212]),.outp(outp[239:160])); 

dbram_4096_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[423:318]),.outp(outp[319:240])); 

dbram_4096_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[529:424]),.outp(outp[399:320])); 

dbram_4096_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[635:530]),.outp(outp[479:400])); 

dbram_4096_40bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[741:636]),.outp(outp[559:480])); 

dbram_4096_40bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[847:742]),.outp(outp[639:560])); 

dbram_4096_40bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[953:848]),.outp(outp[719:640])); 

dbram_4096_40bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1059:954]),.outp(outp[799:720])); 

endmodule 



module dbram_4096_60bit_module_20(input clk, input reset, input[2919:0] inp, output [2399:0] outp); 

dbram_4096_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[145:0]),.outp(outp[119:0])); 

dbram_4096_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[291:146]),.outp(outp[239:120])); 

dbram_4096_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[437:292]),.outp(outp[359:240])); 

dbram_4096_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[583:438]),.outp(outp[479:360])); 

dbram_4096_60bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[729:584]),.outp(outp[599:480])); 

dbram_4096_60bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[875:730]),.outp(outp[719:600])); 

dbram_4096_60bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1021:876]),.outp(outp[839:720])); 

dbram_4096_60bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[1167:1022]),.outp(outp[959:840])); 

dbram_4096_60bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[1313:1168]),.outp(outp[1079:960])); 

dbram_4096_60bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1459:1314]),.outp(outp[1199:1080])); 

dbram_4096_60bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[1605:1460]),.outp(outp[1319:1200])); 

dbram_4096_60bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[1751:1606]),.outp(outp[1439:1320])); 

dbram_4096_60bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[1897:1752]),.outp(outp[1559:1440])); 

dbram_4096_60bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[2043:1898]),.outp(outp[1679:1560])); 

dbram_4096_60bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[2189:2044]),.outp(outp[1799:1680])); 

dbram_4096_60bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[2335:2190]),.outp(outp[1919:1800])); 

dbram_4096_60bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[2481:2336]),.outp(outp[2039:1920])); 

dbram_4096_60bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[2627:2482]),.outp(outp[2159:2040])); 

dbram_4096_60bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[2773:2628]),.outp(outp[2279:2160])); 

dbram_4096_60bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[2919:2774]),.outp(outp[2399:2280])); 

endmodule 

module activation_32_16bit_module_6(input clk, input reset, input[3095:0] inp, output [3083:0] outp); 

activation_32_16bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[515:0]),.outp(outp[513:0])); 

activation_32_16bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[1031:516]),.outp(outp[1027:514])); 

activation_32_16bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[1547:1032]),.outp(outp[1541:1028])); 

activation_32_16bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[2063:1548]),.outp(outp[2055:1542])); 

activation_32_16bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[2579:2064]),.outp(outp[2569:2056])); 

activation_32_16bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[3095:2580]),.outp(outp[3083:2570])); 

endmodule 

module activation_32_8bit_module_12(input clk, input reset, input[3131:0] inp, output [3095:0] outp); 

activation_32_8bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[260:0]),.outp(outp[257:0])); 

activation_32_8bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[521:261]),.outp(outp[515:258])); 

activation_32_8bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[782:522]),.outp(outp[773:516])); 

activation_32_8bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1043:783]),.outp(outp[1031:774])); 

activation_32_8bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[1304:1044]),.outp(outp[1289:1032])); 

activation_32_8bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1565:1305]),.outp(outp[1547:1290])); 

activation_32_8bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1826:1566]),.outp(outp[1805:1548])); 

activation_32_8bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[2087:1827]),.outp(outp[2063:1806])); 

activation_32_8bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[2348:2088]),.outp(outp[2321:2064])); 

activation_32_8bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[2609:2349]),.outp(outp[2579:2322])); 

activation_32_8bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[2870:2610]),.outp(outp[2837:2580])); 

activation_32_8bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[3131:2871]),.outp(outp[3095:2838])); 

endmodule 

module adder_tree_3_8bit_14(input clk, input reset, input[895:0] inp, output [223:0] outp); 

adder_tree_3_8bit inst_0 (.clk(clk),.reset(reset),.inp(inp[63:0]),.outp(outp[15:0])); 

adder_tree_3_8bit inst_1 (.clk(clk),.reset(reset),.inp(inp[127:64]),.outp(outp[31:16])); 

adder_tree_3_8bit inst_2 (.clk(clk),.reset(reset),.inp(inp[191:128]),.outp(outp[47:32])); 

adder_tree_3_8bit inst_3 (.clk(clk),.reset(reset),.inp(inp[255:192]),.outp(outp[63:48])); 

adder_tree_3_8bit inst_4 (.clk(clk),.reset(reset),.inp(inp[319:256]),.outp(outp[79:64])); 

adder_tree_3_8bit inst_5 (.clk(clk),.reset(reset),.inp(inp[383:320]),.outp(outp[95:80])); 

adder_tree_3_8bit inst_6 (.clk(clk),.reset(reset),.inp(inp[447:384]),.outp(outp[111:96])); 

adder_tree_3_8bit inst_7 (.clk(clk),.reset(reset),.inp(inp[511:448]),.outp(outp[127:112])); 

adder_tree_3_8bit inst_8 (.clk(clk),.reset(reset),.inp(inp[575:512]),.outp(outp[143:128])); 

adder_tree_3_8bit inst_9 (.clk(clk),.reset(reset),.inp(inp[639:576]),.outp(outp[159:144])); 

adder_tree_3_8bit inst_10 (.clk(clk),.reset(reset),.inp(inp[703:640]),.outp(outp[175:160])); 

adder_tree_3_8bit inst_11 (.clk(clk),.reset(reset),.inp(inp[767:704]),.outp(outp[191:176])); 

adder_tree_3_8bit inst_12 (.clk(clk),.reset(reset),.inp(inp[831:768]),.outp(outp[207:192])); 

adder_tree_3_8bit inst_13 (.clk(clk),.reset(reset),.inp(inp[895:832]),.outp(outp[223:208])); 

endmodule 

module adder_tree_4_4bit_24(input clk, input reset, input[1535:0] inp, output [191:0] outp); 

adder_tree_4_4bit inst_0 (.clk(clk),.reset(reset),.inp(inp[63:0]),.outp(outp[7:0])); 

adder_tree_4_4bit inst_1 (.clk(clk),.reset(reset),.inp(inp[127:64]),.outp(outp[15:8])); 

adder_tree_4_4bit inst_2 (.clk(clk),.reset(reset),.inp(inp[191:128]),.outp(outp[23:16])); 

adder_tree_4_4bit inst_3 (.clk(clk),.reset(reset),.inp(inp[255:192]),.outp(outp[31:24])); 

adder_tree_4_4bit inst_4 (.clk(clk),.reset(reset),.inp(inp[319:256]),.outp(outp[39:32])); 

adder_tree_4_4bit inst_5 (.clk(clk),.reset(reset),.inp(inp[383:320]),.outp(outp[47:40])); 

adder_tree_4_4bit inst_6 (.clk(clk),.reset(reset),.inp(inp[447:384]),.outp(outp[55:48])); 

adder_tree_4_4bit inst_7 (.clk(clk),.reset(reset),.inp(inp[511:448]),.outp(outp[63:56])); 

adder_tree_4_4bit inst_8 (.clk(clk),.reset(reset),.inp(inp[575:512]),.outp(outp[71:64])); 

adder_tree_4_4bit inst_9 (.clk(clk),.reset(reset),.inp(inp[639:576]),.outp(outp[79:72])); 

adder_tree_4_4bit inst_10 (.clk(clk),.reset(reset),.inp(inp[703:640]),.outp(outp[87:80])); 

adder_tree_4_4bit inst_11 (.clk(clk),.reset(reset),.inp(inp[767:704]),.outp(outp[95:88])); 

adder_tree_4_4bit inst_12 (.clk(clk),.reset(reset),.inp(inp[831:768]),.outp(outp[103:96])); 

adder_tree_4_4bit inst_13 (.clk(clk),.reset(reset),.inp(inp[895:832]),.outp(outp[111:104])); 

adder_tree_4_4bit inst_14 (.clk(clk),.reset(reset),.inp(inp[959:896]),.outp(outp[119:112])); 

adder_tree_4_4bit inst_15 (.clk(clk),.reset(reset),.inp(inp[1023:960]),.outp(outp[127:120])); 

adder_tree_4_4bit inst_16 (.clk(clk),.reset(reset),.inp(inp[1087:1024]),.outp(outp[135:128])); 

adder_tree_4_4bit inst_17 (.clk(clk),.reset(reset),.inp(inp[1151:1088]),.outp(outp[143:136])); 

adder_tree_4_4bit inst_18 (.clk(clk),.reset(reset),.inp(inp[1215:1152]),.outp(outp[151:144])); 

adder_tree_4_4bit inst_19 (.clk(clk),.reset(reset),.inp(inp[1279:1216]),.outp(outp[159:152])); 

adder_tree_4_4bit inst_20 (.clk(clk),.reset(reset),.inp(inp[1343:1280]),.outp(outp[167:160])); 

adder_tree_4_4bit inst_21 (.clk(clk),.reset(reset),.inp(inp[1407:1344]),.outp(outp[175:168])); 

adder_tree_4_4bit inst_22 (.clk(clk),.reset(reset),.inp(inp[1471:1408]),.outp(outp[183:176])); 

adder_tree_4_4bit inst_23 (.clk(clk),.reset(reset),.inp(inp[1535:1472]),.outp(outp[191:184])); 

endmodule 

module adder_tree_4_16bit_20(input clk, input reset, input[5119:0] inp, output [639:0] outp); 

adder_tree_4_16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[255:0]),.outp(outp[31:0])); 

adder_tree_4_16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[511:256]),.outp(outp[63:32])); 

adder_tree_4_16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[767:512]),.outp(outp[95:64])); 

adder_tree_4_16bit inst_3 (.clk(clk),.reset(reset),.inp(inp[1023:768]),.outp(outp[127:96])); 

adder_tree_4_16bit inst_4 (.clk(clk),.reset(reset),.inp(inp[1279:1024]),.outp(outp[159:128])); 

adder_tree_4_16bit inst_5 (.clk(clk),.reset(reset),.inp(inp[1535:1280]),.outp(outp[191:160])); 

adder_tree_4_16bit inst_6 (.clk(clk),.reset(reset),.inp(inp[1791:1536]),.outp(outp[223:192])); 

adder_tree_4_16bit inst_7 (.clk(clk),.reset(reset),.inp(inp[2047:1792]),.outp(outp[255:224])); 

adder_tree_4_16bit inst_8 (.clk(clk),.reset(reset),.inp(inp[2303:2048]),.outp(outp[287:256])); 

adder_tree_4_16bit inst_9 (.clk(clk),.reset(reset),.inp(inp[2559:2304]),.outp(outp[319:288])); 

adder_tree_4_16bit inst_10 (.clk(clk),.reset(reset),.inp(inp[2815:2560]),.outp(outp[351:320])); 

adder_tree_4_16bit inst_11 (.clk(clk),.reset(reset),.inp(inp[3071:2816]),.outp(outp[383:352])); 

adder_tree_4_16bit inst_12 (.clk(clk),.reset(reset),.inp(inp[3327:3072]),.outp(outp[415:384])); 

adder_tree_4_16bit inst_13 (.clk(clk),.reset(reset),.inp(inp[3583:3328]),.outp(outp[447:416])); 

adder_tree_4_16bit inst_14 (.clk(clk),.reset(reset),.inp(inp[3839:3584]),.outp(outp[479:448])); 

adder_tree_4_16bit inst_15 (.clk(clk),.reset(reset),.inp(inp[4095:3840]),.outp(outp[511:480])); 

adder_tree_4_16bit inst_16 (.clk(clk),.reset(reset),.inp(inp[4351:4096]),.outp(outp[543:512])); 

adder_tree_4_16bit inst_17 (.clk(clk),.reset(reset),.inp(inp[4607:4352]),.outp(outp[575:544])); 

adder_tree_4_16bit inst_18 (.clk(clk),.reset(reset),.inp(inp[4863:4608]),.outp(outp[607:576])); 

adder_tree_4_16bit inst_19 (.clk(clk),.reset(reset),.inp(inp[5119:4864]),.outp(outp[639:608])); 

endmodule 


module dbram_2048_60bit_module_1(input clk, input reset, input[143:0] inp, output [119:0] outp); 

dbram_2048_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[143:0]),.outp(outp[119:0])); 

endmodule 

module systolic_array_4_fp16bit_1(input clk, input reset, input[417:0] inp, output [223:0] outp); 

systolic_array_4_fp16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[417:0]),.outp(outp[223:0])); 

endmodule 

module sigmoid_16bit_8(input clk, input reset, input[127:0] inp, output [127:0] outp); 

sigmoid_16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[15:0]),.outp(outp[15:0])); 

sigmoid_16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[31:16]),.outp(outp[31:16])); 

sigmoid_16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[47:32]),.outp(outp[47:32])); 

sigmoid_16bit inst_3 (.clk(clk),.reset(reset),.inp(inp[63:48]),.outp(outp[63:48])); 

sigmoid_16bit inst_4 (.clk(clk),.reset(reset),.inp(inp[79:64]),.outp(outp[79:64])); 

sigmoid_16bit inst_5 (.clk(clk),.reset(reset),.inp(inp[95:80]),.outp(outp[95:80])); 

sigmoid_16bit inst_6 (.clk(clk),.reset(reset),.inp(inp[111:96]),.outp(outp[111:96])); 

sigmoid_16bit inst_7 (.clk(clk),.reset(reset),.inp(inp[127:112]),.outp(outp[127:112])); 

endmodule 

module adder_tree_3_8bit_6(input clk, input reset, input[383:0] inp, output [95:0] outp); 

adder_tree_3_8bit inst_0 (.clk(clk),.reset(reset),.inp(inp[63:0]),.outp(outp[15:0])); 

adder_tree_3_8bit inst_1 (.clk(clk),.reset(reset),.inp(inp[127:64]),.outp(outp[31:16])); 

adder_tree_3_8bit inst_2 (.clk(clk),.reset(reset),.inp(inp[191:128]),.outp(outp[47:32])); 

adder_tree_3_8bit inst_3 (.clk(clk),.reset(reset),.inp(inp[255:192]),.outp(outp[63:48])); 

adder_tree_3_8bit inst_4 (.clk(clk),.reset(reset),.inp(inp[319:256]),.outp(outp[79:64])); 

adder_tree_3_8bit inst_5 (.clk(clk),.reset(reset),.inp(inp[383:320]),.outp(outp[95:80])); 

endmodule 

module adder_tree_4_4bit_18(input clk, input reset, input[1151:0] inp, output [143:0] outp); 

adder_tree_4_4bit inst_0 (.clk(clk),.reset(reset),.inp(inp[63:0]),.outp(outp[7:0])); 

adder_tree_4_4bit inst_1 (.clk(clk),.reset(reset),.inp(inp[127:64]),.outp(outp[15:8])); 

adder_tree_4_4bit inst_2 (.clk(clk),.reset(reset),.inp(inp[191:128]),.outp(outp[23:16])); 

adder_tree_4_4bit inst_3 (.clk(clk),.reset(reset),.inp(inp[255:192]),.outp(outp[31:24])); 

adder_tree_4_4bit inst_4 (.clk(clk),.reset(reset),.inp(inp[319:256]),.outp(outp[39:32])); 

adder_tree_4_4bit inst_5 (.clk(clk),.reset(reset),.inp(inp[383:320]),.outp(outp[47:40])); 

adder_tree_4_4bit inst_6 (.clk(clk),.reset(reset),.inp(inp[447:384]),.outp(outp[55:48])); 

adder_tree_4_4bit inst_7 (.clk(clk),.reset(reset),.inp(inp[511:448]),.outp(outp[63:56])); 

adder_tree_4_4bit inst_8 (.clk(clk),.reset(reset),.inp(inp[575:512]),.outp(outp[71:64])); 

adder_tree_4_4bit inst_9 (.clk(clk),.reset(reset),.inp(inp[639:576]),.outp(outp[79:72])); 

adder_tree_4_4bit inst_10 (.clk(clk),.reset(reset),.inp(inp[703:640]),.outp(outp[87:80])); 

adder_tree_4_4bit inst_11 (.clk(clk),.reset(reset),.inp(inp[767:704]),.outp(outp[95:88])); 

adder_tree_4_4bit inst_12 (.clk(clk),.reset(reset),.inp(inp[831:768]),.outp(outp[103:96])); 

adder_tree_4_4bit inst_13 (.clk(clk),.reset(reset),.inp(inp[895:832]),.outp(outp[111:104])); 

adder_tree_4_4bit inst_14 (.clk(clk),.reset(reset),.inp(inp[959:896]),.outp(outp[119:112])); 

adder_tree_4_4bit inst_15 (.clk(clk),.reset(reset),.inp(inp[1023:960]),.outp(outp[127:120])); 

adder_tree_4_4bit inst_16 (.clk(clk),.reset(reset),.inp(inp[1087:1024]),.outp(outp[135:128])); 

adder_tree_4_4bit inst_17 (.clk(clk),.reset(reset),.inp(inp[1151:1088]),.outp(outp[143:136])); 

endmodule 
module adder_tree_1_16bit (input clk,input reset,input [31:0] inp, output [31:0] outp);

adder_tree_1stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.sum_out(outp));

endmodule

module adder_tree_2_16bit (input clk, input reset, input [63:0] inp, output [31:0] outp);

adder_tree_2stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.sum_out(outp));

endmodule

module adder_tree_3_16bit (input clk, input reset, input [127:0] inp, output [31:0] outp);

adder_tree_3stage_16bit inst (.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.inp20(inp[79:64]),.inp21(inp[95:80]),.inp30(inp[111:96]),.inp31(inp[127:112]),.sum_out(outp));

endmodule

module adder_tree_4_16bit (input clk, input reset, input [255:0] inp, output [31:0] outp);

adder_tree_4stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.inp20(inp[79:64]),.inp21(inp[95:80]),.inp30(inp[111:96]),.inp31(inp[127:112]),.inp40(inp[143:128]),.inp41(inp[159:144]),.inp50(inp[175:160]),.inp51(inp[191:176]),.inp60(inp[207:192]),.inp61(inp[223:208]),.inp70(inp[239:224]),.inp71(inp[255:240]),.sum_out(outp));

endmodule

module adder_tree_1_8bit (input clk, input reset, input [15:0] inp, output [15:0] outp);

adder_tree_1stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.sum_out(outp));

endmodule

module adder_tree_2_8bit (input clk, input reset, input [31:0] inp, output [15:0] outp);

adder_tree_2stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.sum_out(outp));

endmodule

module adder_tree_3_8bit (input clk, input reset, input [63:0] inp, output [15:0] outp);

adder_tree_3stage_8bit inst (.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.inp20(inp[39:32]),.inp21(inp[47:40]),.inp30(inp[55:48]),.inp31(inp[63:56]),.sum_out(outp));

endmodule

module adder_tree_4_8bit (input clk, input reset, input [127:0] inp, output [15:0] outp);

adder_tree_4stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.inp20(inp[39:32]),.inp21(inp[47:40]),.inp30(inp[55:48]),.inp31(inp[63:56]),.inp40(inp[71:64]),.inp41(inp[79:72]),.inp50(inp[87:80]),.inp51(inp[95:88]),.inp60(inp[103:96]),.inp61(inp[111:104]),.inp70(inp[119:112]),.inp71(inp[127:120]),.sum_out(outp));

endmodule

module adder_tree_1_4bit (input clk, input reset, input [7:0] inp, output [7:0] outp);

adder_tree_1stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.sum_out(outp));

endmodule

module adder_tree_2_4bit (input clk, input reset, input [15:0] inp, output [7:0] outp);

adder_tree_2stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.sum_out(outp));

endmodule

module adder_tree_3_4bit (input clk, input reset, input [31:0] inp, output [7:0] outp);

adder_tree_3stage_4bit inst (.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.inp20(inp[19:16]),.inp21(inp[23:20]),.inp30(inp[27:24]),.inp31(inp[31:28]),.sum_out(outp));

endmodule

module adder_tree_4_4bit (input clk, input reset, input [63:0] inp, output [7:0] outp);

adder_tree_4stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.inp20(inp[19:16]),.inp21(inp[23:20]),.inp30(inp[27:24]),.inp31(inp[31:28]),.inp40(inp[35:32]),.inp41(inp[39:36]),.inp50(inp[43:40]),.inp51(inp[47:44]),.inp60(inp[51:48]),.inp61(inp[55:52]),.inp70(inp[59:56]),.inp71(inp[63:60]),.sum_out(outp));

endmodule

module adder_tree_3_fp16bit (input clk, input reset, input [131:0] inp, output [15:0] outp);

mode4_adder_tree inst(
  .inp0(inp[15:0]),
  .inp1(inp[31:16]),
  .inp2(inp[47:32]),
  .inp3(inp[63:48]),
  .inp4(inp[79:64]),
  .inp5(inp[95:80]),
  .inp6(inp[111:96]),
  .inp7(inp[127:112]),
  .mode4_stage0_run(inp[128]),
  .mode4_stage1_run(inp[129]),
  .mode4_stage2_run(inp[130]),
  .mode4_stage3_run(inp[131]),

  .clk(clk),
  .reset(reset),
  .outp(outp[15:0])
);

endmodule

module dpram_1024_32bit_module (input clk, input reset, input [85:0] inp, output [63:0] outp);

dpram inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[53:22]),.data_b(inp[85:54]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_1024_64bit_module (input clk, input reset, input [149:0] inp, output [63:0] outp );

dpram_1024_64bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[85:22]),.data_b(inp[149:86]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_2048_64bit_module (input clk, input reset, input [151:0] inp, output [127:0] outp);

dpram_2048_64bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[87:24]),.data_b(inp[151:88]),.out_a(outp[63:0]),.out_b(outp[127:64]));

endmodule

module dpram_2048_32bit_module (input clk, input reset, input [87:0] inp, output [63:0] outp);

dpram_2048_32bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[55:24]),.data_b(inp[87:56]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_1024_40bit_module (input clk, input reset, input [101:0] inp, output [79:0] outp);

dpram_1024_40bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[61:22]),.data_b(inp[101:62]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_1024_60bit_module (input clk, input reset, input [141:0] inp, output [119:0] outp);

dpram_1024_60bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[81:22]),.data_b(inp[141:82]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dpram_2048_40bit_module (input clk, input reset, input [103:0] inp, output [79:0] outp);

dpram_2048_40bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[63:24]),.data_b(inp[103:64]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_2048_60bit_module (input clk, input reset, input [143:0] inp, output [119:0] outp);

dpram_2048_60bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[83:24]),.data_b(inp[143:84]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dpram_4096_40bit_module (input clk, input reset, input [105:0] inp, output [79:0] outp);

dpram_4096_40bit inst (.clk(clk),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[65:26]),.data_b(inp[105:66]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_4096_60bit_module (input clk, input reset, input [145:0] inp, output [119:0] outp);

dpram_4096_60bit inst (.clk(clk),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[85:26]),.data_b(inp[145:86]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module spram_1024_32bit_module (input clk,input reset,input [42:0] inp, output [31:0] outp);

spram inst (.clk(clk),.address(inp[9:0]),.wren(inp[10]),.data(inp[42:11]),.out(outp));

endmodule

module spram_2048_40bit_module (input clk,input reset,input [51:0] inp, output [39:0] outp);

spram_2048_40bit inst (.clk(clk),.address(inp[10:0]),.wren(inp[11]),.data(inp[51:12]),.out(outp));

endmodule

module spram_2048_60bit_module (input clk,input reset,input [71:0] inp, output [59:0] outp);

spram_2048_60bit inst (.clk(clk),.address(inp[10:0]),.wren(inp[11]),.data(inp[71:12]),.out(outp));

endmodule

module spram_4096_40bit_module (input clk,input reset,input [52:0] inp, output [39:0] outp);

spram_4096_40bit inst (.clk(clk),.address(inp[11:0]),.wren(inp[12]),.data(inp[52:13]),.out(outp));

endmodule

module spram_4096_60bit_module (input clk,input reset,input [72:0] inp, output [59:0] outp);

spram_4096_60bit inst (.clk(clk),.address(inp[11:0]),.wren(inp[12]),.data(inp[72:13]),.out(outp));

endmodule

module dbram_2048_40bit_module (input clk,input reset,input [103:0] inp, output [79:0] outp);

dbram_2048_40bit inst (.clk(clk),.reset(reset),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[63:24]),.data_b(inp[103:64]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dbram_2048_60bit_module (input clk,input reset,input [143:0] inp, output [119:0] outp);

dbram_2048_60bit inst (.clk(clk),.reset(reset),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[83:24]),.data_b(inp[143:84]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dbram_4096_40bit_module (input clk,input reset,input [105:0] inp, output [79:0] outp);

dbram_4096_40bit inst (.clk(clk),.reset(reset),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[65:26]),.data_b(inp[105:66]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dbram_4096_60bit_module (input clk,input reset,input [145:0] inp, output [119:0] outp);

dbram_4096_60bit inst (.clk(clk),.reset(reset),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[85:26]),.data_b(inp[145:86]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule


module fifo_256_40bit_module (input clk,input reset,input [42:0] inp, output [41:0] outp);

fifo_256_40bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[40:1]),.we(inp[41]),.dout(outp[39:0]),.re(inp[42]),.full(outp[40]),.empty(outp[41]));

endmodule

module fifo_256_60bit_module (input clk,input reset,input [62:0] inp, output [61:0] outp);

fifo_256_60bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[60:1]),.we(inp[61]),.dout(outp[59:0]),.re(inp[62]),.full(outp[60]),.empty(outp[61]));

endmodule

module fifo_512_60bit_module (input clk,input reset,input [62:0] inp, output [61:0] outp);

fifo_512_60bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[60:1]),.we(inp[61]),.dout(outp[59:0]),.re(inp[62]),.full(outp[60]),.empty(outp[61]));

endmodule

module fifo_512_40bit_module (input clk,input reset,input [42:0] inp, output [41:0] outp);

fifo_512_40bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[40:1]),.we(inp[41]),.dout(outp[39:0]),.re(inp[42]),.full(outp[40]),.empty(outp[41]));

endmodule

module tanh_16bit (input clk,input reset, input [15:0] inp, output [15:0] outp);

tanh inst (.x(inp),.tanh_out(outp));

endmodule

module sigmoid_16bit (input clk,input reset, input [15:0] inp, output [15:0] outp);

sigmoid inst (.x(inp),.sig_out(outp));

endmodule

module systolic_array_4_16bit (input clk, input reset, input [254:0] inp, output [130:0] outp);

matmul_4x4_systolic inst(
 .clk(clk),
 .reset(inp[254]),
 .pe_reset(reset),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[11:1]),
 .address_mat_b(inp[22:12]),
 .address_mat_c(inp[33:23]),
 .address_stride_a(inp[41:34]),
 .address_stride_b(inp[49:42]),
 .address_stride_c(inp[57:50]),
 .a_data(inp[89:58]),
 .b_data(inp[121:90]),
 .a_data_in(inp[153:122]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[185:154]),
 .c_data_in(inp[217:186]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[32:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[64:33]),
 .b_data_out(outp[96:65]),
 .a_addr(outp[107:97]),
 .b_addr(outp[118:108]),
 .c_addr(outp[129:119]),
 .c_data_available(outp[130]),
 .validity_mask_a_rows(inp[221:218]),
 .validity_mask_a_cols_b_rows(inp[225:222]),
 .validity_mask_b_cols(inp[229:226]),
 .final_mat_mul_size(inp[237:230]),
 .a_loc(inp[245:238]),
 .b_loc(inp[253:246])
);

endmodule

module systolic_array_8_16bit (input clk, input reset, input [785:0] inp, output [433:0] outp);

matmul_8x8_systolic inst(
 .clk(clk),
 .reset(reset),
 .pe_reset(inp[785]),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[16:1]),
 .address_mat_b(inp[32:17]),
 .address_mat_c(inp[48:33]),
 .address_stride_a(inp[64:49]),
 .address_stride_b(inp[80:65]),
 .address_stride_c(inp[96:81]),
 .a_data(inp[224:97]),
 .b_data(inp[352:225]),
 .a_data_in(inp[480:353]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[608:481]),
 .c_data_in(inp[736:609]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[128:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[256:129]),
 .b_data_out(outp[384:257]),
 .a_addr(outp[400:385]),
 .b_addr(outp[416:401]),
 .c_addr(outp[432:417]),
 .c_data_available(outp[433]),
 .validity_mask_a_rows(inp[744:737]),
 .validity_mask_a_cols_b_rows(inp[752:745]),
 .validity_mask_b_cols(inp[760:753]),
 .final_mat_mul_size(inp[768:761]),
 .a_loc(inp[776:769]),
 .b_loc(inp[784:777])
);

endmodule

module systolic_array_4_fp16bit (input clk, input reset, input [417:0] inp, output [223:0] outp);

matmul_4x4_fp_systolic inst(
 .clk(clk),
 .reset(reset),
 .pe_reset(inp[417]),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[10:1]),
 .address_mat_b(inp[20:11]),
 .address_mat_c(inp[30:21]),
 .address_stride_a(inp[40:31]),
 .address_stride_b(inp[50:41]),
 .address_stride_c(inp[60:51]),
 .a_data(inp[124:61]),
 .b_data(inp[188:125]),
 .a_data_in(inp[252:189]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[316:253]),
 .c_data_in(inp[380:317]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[64:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[128:65]),
 .b_data_out(outp[192:129]),
 .a_addr(outp[202:193]),
 .b_addr(outp[212:203]),
 .c_addr(outp[222:213]),
 .c_data_available(outp[223]),
 .validity_mask_a_rows(inp[384:381]),
 .validity_mask_a_cols_b_rows(inp[388:385]),
 .validity_mask_b_cols(inp[392:389]),
 .final_mat_mul_size(inp[400:393]),
 .a_loc(inp[408:401]),
 .b_loc(inp[416:409])
);

endmodule

module dsp_chain_2_int_sop_2_module (input clk, input reset, input [147:0] inp, output [36:0] outp);

dsp_chain_2_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.result(outp[36:0]));

endmodule

module dsp_chain_3_int_sop_2_module (input clk, input reset, input [221:0] inp, output [36:0] outp);

dsp_chain_3_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.ax3(inp[165:148]),.ay3(inp[184:166]),.bx3(inp[202:185]),.by3(inp[221:203]),.result(outp[36:0]));

endmodule

module dsp_chain_4_int_sop_2_module (input clk, input reset, input [295:0] inp, output [36:0] outp);

dsp_chain_4_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.ax3(inp[165:148]),.ay3(inp[184:166]),.bx3(inp[202:185]),.by3(inp[221:203]),.ax4(inp[239:222]),.ay4(inp[258:240]),.bx4(inp[276:259]),.by4(inp[295:277]),.result(outp[36:0]));

endmodule

module dsp_chain_2_fp16_sop2_mult_module (input clk, input reset, input [127:0] inp, output [31:0] outp);

dsp_chain_2_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.result(outp));

endmodule

module dsp_chain_3_fp16_sop2_mult_module (input clk, input reset, input [191:0] inp, output [31:0] outp);

dsp_chain_3_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.top_a3(inp[143:128]),.top_b3(inp[159:144]),.bot_a3(inp[175:160]),.bot_b3(inp[191:176]),.result(outp));

endmodule

module dsp_chain_4_fp16_sop2_mult_module (input clk, input reset, input [255:0] inp, output [31:0] outp);

dsp_chain_4_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.top_a3(inp[143:128]),.top_b3(inp[159:144]),.bot_a3(inp[175:160]),.bot_b3(inp[191:176]),.top_a4(inp[207:192]),.top_b4(inp[223:208]),.bot_a4(inp[239:224]),.bot_b4(inp[255:240]),.result(outp));

endmodule

module tensor_block_bf16_module (input clk, input reset, input [264:0] inp, output [271:0] outp);

tensor_block_bf16 inst(
	.clk(clk),
	.reset(reset),

	.data_in(inp[79:0]),
	.cascade_in(inp[159:80]),
	.acc0_in(inp[191:160]),
	.acc1_in(inp[223:192]),
	.acc2_in(inp[255:224]),
	.accumulator_input1_select(inp[258:256]),

	.out0(outp[31:0]),
	.out1(outp[63:32]),
	.out2(outp[95:64]),
	.cascade_out(outp[175:96]),
	.acc0_out(outp[207:176]),
	.acc1_out(outp[239:208]),
	.acc2_out(outp[271:240]),

	.mux1_select(inp[259]),
	.dot_unit_input_1_enable(inp[260]),
	.bank0_data_in_enable(inp[261]),
	.bank1_data_in_enable(inp[262]),
	.cascade_out_select(inp[263]),
	.dot_unit_input_2_select(inp[264])

	);

endmodule

module tensor_block_int8_module (input clk, input reset, input [264:0] inp, output [250:0] outp);

tensor_block inst(
	.clk(clk),
	.reset(reset),

	.data_in(inp[79:0]),
	.cascade_in(inp[159:80]),
	.acc0_in(inp[191:160]),
	.acc1_in(inp[223:192]),
	.acc2_in(inp[255:224]),
	.accumulator_input1_select(inp[258:256]),

	.out0(outp[24:0]),
	.out1(outp[49:25]),
	.out2(outp[74:50]),
	.cascade_out(outp[154:75]),
	.acc0_out(outp[186:155]),
	.acc1_out(outp[218:187]),
	.acc2_out(outp[250:219]),

	.mux1_select(inp[259]),
	.dot_unit_input_1_enable(inp[260]),
	.bank0_data_in_enable(inp[261]),
	.bank1_data_in_enable(inp[262]),
	.cascade_out_select(inp[263]),
	.dot_unit_input_2_select(inp[264])

	);

endmodule


module activation_32_8bit_module (input clk, input reset, input [260:0] inp, output [257:0] outp);

activation_32_8bit inst (
    .activation_type(inp[0]),
    .enable_activation(inp[1]),
    .in_data_available(inp[2]),
    .inp_data(inp[258:3]),
    .out_data(outp[255:0]),
    .out_data_available(outp[256]),
    .validity_mask(inp[260:259]),
    .done_activation(outp[257]),
    .clk(clk),
    .reset(reset)
);

endmodule

module activation_32_16bit_module (input clk, input reset, input [515:0] inp, output [513:0] outp);

activation_32_16bit inst (
    .activation_type(inp[0]),
    .enable_activation(inp[1]),
    .in_data_available(inp[2]),
    .inp_data(inp[514:3]),
    .out_data(outp[511:0]),
    .out_data_available(outp[512]),
    .validity_mask(inp[515:514]),
    .done_activation(outp[513]),
    .clk(clk),
    .reset(reset)
);

endmodule

module fsm(input clk, input reset, input i1, input i2, output reg o);
// mealy machine

reg [1:0] current_state; 
reg [1:0] next_state;

wire [1:0] inp; 
assign inp = {i2,i1}; 

always@(posedge clk) begin 
	if (reset == 1'b1) begin 
		current_state <= 1'b0; 
	end
	else begin 
		current_state <= next_state; 
	end
end

always@(posedge clk) begin 

	next_state = current_state; 

	case(current_state)
		2'b00:	begin 
							if(inp == 2'b00) begin 
								next_state <= 2'b00; 
								o <= 1'b0; 
							end
							if (inp == 2'b01) begin 
								next_state <= 2'b11;
								o <= 1'b1;
							end
							if(inp == 2'b10) begin
  							next_state <= 2'b01;
  							o <= 1'b0;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b10;
							  o <= 1'b0;
							end
					 	end 
		2'b01:	begin 
							if(inp == 2'b00) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b01;
							  o <= 1'b0;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b00;
							  o <= 1'b1;
							end
						end
		2'b10:	begin 
							if(inp == 2'b00) begin
							  next_state <= 2'b11;
							  o <= 1'b0;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b11;
							  o <= 1'b0;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
						end
		2'b11:	begin 
							if(inp == 2'b00) begin
  							next_state <= 2'b00;
							  o <= 1'b1;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b11;
							  o <= 1'b1;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
						end
//		defualt:	begin  
//								next_state <= 2'b00;
//								o <= 1'b0; 
//							end
	endcase
end 

endmodule 
module xor_module (input clk, input reset, input i1, input i2, output reg o);

always@(posedge clk) begin 
if (reset ==1'b1) begin 
o<= 1'b0; 
end
else begin
o <= i1^i2; 
end 
end
endmodule
module mux_module (input clk, input reset, input i1, input i2, output reg o, input sel);

always@(posedge clk) begin 
if (reset ==1'b1) begin 
	o<= 1'b0; 
end

else begin
	if (sel == 1'b0) begin 
		o <= i1;
	end
	else begin
		o <= i2; 
	end 
end 

end

endmodule

`ifdef complex_dsp
module int_sop_2_dspchain (mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
	chainin,
	resulta,
	chainout);
input [10:0] mode_sigs;
input clk;
input reset; 
input [17:0] ax, bx;
input [18:0] ay, by;
input [36:0] chainin;

output [36:0] resulta;
output [36:0] chainout;

wire [11:0] mode_sigs_int;
assign mode_sigs_int = {1'b0, mode_sigs};

int_sop_2 inst1(.clk(clk),.reset(reset),.ax(ax),.bx(bx),.ay(ay),.by(by),.mode_sigs(mode_sigs_int),.chainin(chainin),.result(resulta),.chainout(chainout)); 

endmodule
`else
module int_sop_2_dspchain (mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
	chainin,
	resulta,
	chainout);
input [10:0] mode_sigs;
input clk;
input reset; 
input [17:0] ax, bx;
input [18:0] ay, by;
input [36:0] chainin;

output [36:0] resulta;
output [36:0] chainout;
reg [17:0] ax_reg;
reg [18:0] ay_reg;
reg [17:0] bx_reg;
reg [18:0] by_reg;
reg [36:0] resulta_reg;
reg [36:0] resultaxy_reg;
reg [36:0] resultbxy_reg;
always @(posedge clk) begin
  if(reset) begin
    resulta_reg <= 0;
    ax_reg <= 0;
    ay_reg <= 0;
    bx_reg <= 0;
    by_reg <= 0;
  end
  else begin
    ax_reg <= ax;
    ay_reg <= ay;
    bx_reg <= bx;
    by_reg <= by;
    resultaxy_reg <= ax_reg * ay_reg;
    resultbxy_reg <= bx_reg * by_reg;
    resulta_reg <= resultaxy_reg + resultbxy_reg + chainin;
  end
end
assign resulta = resulta_reg;
assign chainout = resulta_reg;
endmodule
`endif

`ifdef complex_dsp
module fp16_sop2_mult_dspchain (clk,reset,top_a,top_b,bot_a,bot_b,fp32_in,mode_sigs,chainin,chainout,result);
input clk; 
input reset;
input [10:0] mode_sigs; 
input [15:0] top_a,top_b,bot_a,bot_b;
input [31:0] chainin,fp32_in; 
output [31:0] chainout, result;

fp16_sop2_mult inst1(.clk(clk),.reset(reset),.top_a(top_a),.top_b(top_b),.bot_a(bot_a),.bot_b(bot_b),.fp32_in(fp32_in),.mode_sigs(mode_sigs),.chainin(chainin),.chainout(chainout),.result(result)); 

endmodule

`else
module fp16_sop2_mult_dspchain (clk,reset,top_a,top_b,bot_a,bot_b,fp32_in,mode_sigs,chainin,chainout,result);
input clk; 
input reset;
input [10:0] mode_sigs; 
input [15:0] top_a,top_b,bot_a,bot_b;
input [31:0] chainin,fp32_in; 
output [31:0] chainout, result; 

reg [15:0] top_a_reg,top_b_reg,bot_a_reg,bot_b_reg; 
reg [31:0] chainin_reg; 
wire [31:0] r1,r2,r3; 
always@(posedge clk) begin 
if(reset) begin 
top_a_reg<= 16'b0; 
top_b_reg<= 16'b0; 
bot_a_reg<= 16'b0; 
bot_b_reg<= 16'b0;
//result<=32'b0;
//chainout<=32'b0;
chainin_reg<=32'b0;   
end
else begin 
top_a_reg<=top_a; 
top_b_reg<=top_b; 
bot_a_reg<=bot_a;
bot_b_reg<=bot_b;
//chainout<=result;
chainin_reg<=chainin; 
end
end

wire [4:0] flags1,flags2,flags3,flags4; 

FPMult_16_dspchain inst1(.clk(clk),.rst(reset),.a(top_a_reg),.b(top_b_reg),.flags(flags1),.result(r1)); 
FPMult_16_dspchain inst2(.clk(clk),.rst(reset),.a(bot_a_reg),.b(bot_b_reg),.flags(flags2),.result(r2));
FPAddSub_single_dspchain inst3(.clk(clk),.rst(reset),.a(r1),.b(r2),.flags(flags3),.operation(1'b1),.result(r3));
FPAddSub_single_dspchain inst4(.clk(clk),.rst(reset),.a(r3),.b(chainin),.flags(flags4),.operation(1'b1),.result(result));
assign chainout = result; 
endmodule
//`endif

//`timescale 1ns / 1ps


// IEEE Half Precision => 5 = 5, 10 = 10



//`define IEEE_COMPLIANCE 1


//////////////////////////////////////////////////////////////////////////////////
//
// Module Name:    FPMult
//
//////////////////////////////////////////////////////////////////////////////////

module FPMult_16_dspchain(
		clk,
		rst,
		a,
		b,
		result,
		flags
    );
	
	// Input Ports
	input clk ;							// Clock
	input rst ;							// Reset signal
	input [16-1:0] a;						// Input A, a 32-bit floating point number
	input [16-1:0] b;						// Input B, a 32-bit floating point number
	
	// Output ports
	output [32-1:0] result ;					// Product, result of the operation, 32-bit FP number
	output [4:0] flags ;						// Flags indicating exceptions according to IEEE754
	
	// Internal signals
	wire [32-1:0] Z_int ;					// Product, result of the operation, 32-bit FP number
	wire [4:0] Flags_int ;						// Flags indicating exceptions according to IEEE754
	
	wire Sa ;							// A's sign
	wire Sb ;							// B's sign
	wire Sp ;							// Product sign
	wire [5-1:0] Ea ;					// A's 5
	wire [5-1:0] Eb ;					// B's 5
	wire [2*10+1:0] Mp ;					// Product 10
	wire [4:0] InputExc ;						// Exceptions in inputs
	wire [23-1:0] NormM ;					// Normalized 10
	wire [8:0] NormE ;					// Normalized 5
	wire [23:0] RoundM ;					// Normalized 10
	wire [8:0] RoundE ;					// Normalized 5
	wire [23:0] RoundMP ;					// Normalized 10
	wire [8:0] RoundEP ;					// Normalized 5
	wire GRS ;

	//reg [63:0] pipe_0;						// Pipeline register Input->Prep
	reg [2*16-1:0] pipe_0;					// Pipeline register Input->Prep

	//reg [92:0] pipe_1;						// Pipeline register Prep->Execute
	//reg [3*10+2*5+7:0] pipe_1;			// Pipeline register Prep->Execute
	reg [3*10+2*5+18:0] pipe_1;

	//reg [38:0] pipe_2;						// Pipeline register Execute->Normalize
	reg [23+8+7:0] pipe_2;				// Pipeline register Execute->Normalize

	//reg [72:0] pipe_3;						// Pipeline register Normalize->Round
	reg [2*23+2*8+10:0] pipe_3;			// Pipeline register Normalize->Round

	//reg [36:0] pipe_4;						// Pipeline register Round->Output
	reg [32+4:0] pipe_4;					// Pipeline register Round->Output
	
	assign result = pipe_4[32+4:5] ;
	assign flags = pipe_4[4:0] ;
	
	// Prepare the operands for alignment and check for exceptions
	FPMult_PrepModule_dspchain PrepModule(clk, rst, pipe_0[2*16-1:16], pipe_0[16-1:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10+1:0], InputExc[4:0]) ;

	// Perform (unsigned) 10 multiplication
	FPMult_ExecuteModule_dspchain ExecuteModule(pipe_1[3*10+5*2+7:2*10+2*5+8], pipe_1[2*10+2*5+7:2*10+7], pipe_1[2*10+6:5], pipe_1[2*10+2*5+6:2*10+5+7], pipe_1[2*10+5+6:2*10+7], pipe_1[2*10+2*5+8], pipe_1[2*10+2*5+7], Sp, NormE[8:0], NormM[23-1:0], GRS) ;

	// Round result and if necessary, perform a second (post-rounding) normalization step
	FPMult_NormalizeModule_dspchain NormalizeModule(pipe_2[23-1:0], pipe_2[23+8:23], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]) ;		

	// Round result and if necessary, perform a second (post-rounding) normalization step
	//FPMult_RoundModule RoundModule(pipe_3[47:24], pipe_3[23:0], pipe_3[65:57], pipe_3[56:48], pipe_3[66], pipe_3[67], pipe_3[72:68], Z_int[31:0], Flags_int[4:0]) ;		
	FPMult_RoundModule_dspchain RoundModule(pipe_3[2*23+1:23+1], pipe_3[23:0], pipe_3[2*8+2*23+3:2*23+8+3], pipe_3[2*23+8+2:2*23+2], pipe_3[2*23+2*8+4], pipe_3[2*23+2*8+5], pipe_3[2*23+2*8+10:2*23+2*8+6], Z_int[32-1:0], Flags_int[4:0]) ;		


//adding always@ (*) instead of posedge clock to make design combinational
	always @ (*) begin	
		if(rst) begin
			pipe_0 = 0;
			pipe_1 = 0;
			pipe_2 = 0; 
			pipe_3 = 0;
			pipe_4 = 0;
		end 
		else begin		
			/* PIPE 0
				[2*16-1:16] A
				[16-1:0] B
			*/
                       pipe_0 = {a, b} ;


			/* PIPE 1
				[2*5+3*10 + 18: 2*5+2*10 + 18] //pipe_0[16+10-1:16] , 10 of A
				[2*5+2*10 + 17 :2*5+2*10 + 9] // pipe_0[8:0]
				[2*5+2*10 + 8] Sa
				[2*5+2*10 + 7] Sb
				[2*5+2*10 + 6:5+2*10+7] Ea
				[5 +2*10+6:2*10+7] Eb
				[2*10+1+5:5] Mp
				[4:0] InputExc
			*/
			//pipe_1 <= {pipe_0[16+10-1:16], pipe_0[10_MUL_SPLIT_LSB-1:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10-1:0], InputExc[4:0]} ;
			pipe_1 = {pipe_0[16+10-1:16], pipe_0[8:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10+1:0], InputExc[4:0]} ;
			
			/* PIPE 2
				[8 + 23 + 7:8 + 23 + 3] InputExc
				[8 + 23 + 2] GRS
				[8 + 23 + 1] Sp
				[8 + 23:23] NormE
				[23-1:0] NormM
			*/
			pipe_2 = {pipe_1[4:0], GRS, Sp, NormE[8:0], NormM[23-1:0]} ;
			/* PIPE 3
				[2*8+2*23+10:2*8+2*23+6] InputExc
				[2*8+2*23+5] GRS
				[2*8+2*23+4] Sp	
				[2*8+2*23+3:8+2*23+3] RoundE
				[8+2*23+2:2*23+2] RoundEP
				[2*23+1:23+1] RoundM
				[23:0] RoundMP
			*/
			pipe_3 = {pipe_2[8 + 23 + 7:8 + 23 + 1], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]} ;
			/* PIPE 4
				[16+4:5] Z
				[4:0] Flags
			*/				
			pipe_4 = {Z_int[32-1:0], Flags_int[4:0]} ;
		end
	end
		
endmodule



module FPMult_PrepModule_dspchain (
		clk,
		rst,
		a,
		b,
		Sa,
		Sb,
		Ea,
		Eb,
		Mp,
		InputExc
	);
	
	// Input ports
	input clk ;
	input rst ;
	input [16-1:0] a ;								// Input A, a 32-bit floating point number
	input [16-1:0] b ;								// Input B, a 32-bit floating point number
	
	// Output ports
	output Sa ;										// A's sign
	output Sb ;										// B's sign
	output [5-1:0] Ea ;								// A's 5
	output [5-1:0] Eb ;								// B's 5
	output [2*10+1:0] Mp ;							// 10 product
	output [4:0] InputExc ;						// Input numbers are exceptions
	
	// Internal signals							// If signal is high...
	wire ANaN ;										// A is a signalling NaN
	wire BNaN ;										// B is a signalling NaN
	wire AInf ;										// A is infinity
	wire BInf ;										// B is infinity
    wire [10-1:0] Ma;
    wire [10-1:0] Mb;
	
	assign ANaN = &(a[16-2:10]) &  |(a[16-2:10]) ;			// All one 5 and not all zero 10 - NaN
	assign BNaN = &(b[16-2:10]) &  |(b[10-1:0]);			// All one 5 and not all zero 10 - NaN
	assign AInf = &(a[16-2:10]) & ~|(a[16-2:10]) ;		// All one 5 and all zero 10 - Infinity
	assign BInf = &(b[16-2:10]) & ~|(b[16-2:10]) ;		// All one 5 and all zero 10 - Infinity
	
	// Check for any exceptions and put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	//assign InputExc = {(ANaN | ANaN | BNaN |BNaN), ANaN, ANaN, BNaN,BNaN} ;
	
	// Take input numbers apart
	assign Sa = a[16-1] ;							// A's sign
	assign Sb = b[16-1] ;							// B's sign
	assign Ea = a[16-2:10];						// Store A's 5 in Ea, unless A is an exception
	assign Eb = b[16-2:10];						// Store B's 5 in Eb, unless B is an exception	
//    assign Ma = a[10_MSB:10_LSB];
  //  assign Mb = b[10_MSB:10_LSB];
	

	// Actual 10 multiplication occurs here
	//assign Mp = ({4'b0001, a[10-1:0]}*{4'b0001, b[10-1:9]}) ;
	assign Mp = ({1'b1,a[10-1:0]}*{1'b1, b[10-1:0]}) ;

	
    //We multiply part of the 10 here
    //Full 10 of A
    //Bits 10_MUL_SPLIT_MSB:10_MUL_SPLIT_LSB of B
   // wire [`ACTUAL_10-1:0] inp_A;
   // wire [`ACTUAL_10-1:0] inp_B;
   // assign inp_A = {1'b1, Ma};
   // assign inp_B = {{(10-(10_MUL_SPLIT_MSB-10_MUL_SPLIT_LSB+1)){1'b0}}, 1'b1, Mb[10_MUL_SPLIT_MSB:10_MUL_SPLIT_LSB]};
   // DW02_mult #(`ACTUAL_10,`ACTUAL_10) u_mult(.A(inp_A), .B(inp_B), .TC(1'b0), .PRODUCT(Mp));
endmodule


module FPMult_ExecuteModule_dspchain(
		a,
		b,
		MpC,
		Ea,
		Eb,
		Sa,
		Sb,
		Sp,
		NormE,
		NormM,
		GRS
    );

	// Input ports
	input [10-1:0] a ;
	input [2*5:0] b ;
	input [2*10+1:0] MpC ;
	input [5-1:0] Ea ;						// A's 5
	input [5-1:0] Eb ;						// B's 5
	input Sa ;								// A's sign
	input Sb ;								// B's sign
	
	// Output ports
	output Sp ;								// Product sign
	output [8:0] NormE ;													// Normalized 5
	output [23-1:0] NormM ;												// Normalized 10
	output GRS ;
	
	wire [2*10+1:0] Mp ;
	
	assign Sp = (Sa ^ Sb) ;												// Equal signs give a positive product
	
   // wire [`ACTUAL_10-1:0] inp_a;
   // wire [`ACTUAL_10-1:0] inp_b;
   // assign inp_a = {1'b1, a};
   // assign inp_b = {{(10-10_MUL_SPLIT_LSB){1'b0}}, 1'b0, b};
   // DW02_mult #(`ACTUAL_10,`ACTUAL_10) u_mult(.A(inp_a), .B(inp_b), .TC(1'b0), .PRODUCT(Mp_temp));
   // DW01_add #(2*`ACTUAL_10) u_add(.A(Mp_temp), .B(MpC<<10_MUL_SPLIT_LSB), .CI(1'b0), .SUM(Mp), .CO());

	//assign Mp = (MpC<<(2*5+1)) + ({4'b0001, a[10-1:0]}*{1'b0, b[2*5:0]}) ;
	assign Mp = MpC;


	assign NormM = (Mp[2*10+1] ? Mp[2*10:0] : Mp[2*10-1:0]); 	// Check for overflow
	assign NormE = (Ea + Eb + Mp[2*10+1]);								// If so, increment 5
	
	assign GRS = ((Mp[10]&(Mp[10+1]))|(|Mp[10-1:0])) ;
	
endmodule

module FPMult_NormalizeModule_dspchain(
		NormM,
		NormE,
		RoundE,
		RoundEP,
		RoundM,
		RoundMP
    );

	// Input Ports
	input [23-1:0] NormM ;									// Normalized 10
	input [8:0] NormE ;									// Normalized 5

	// Output Ports
	output [8:0] RoundE ;
	output [8:0] RoundEP ;
	output [23:0] RoundM ;
	output [23:0] RoundMP ; 
	
// 5 = 5 
// 5 -1 = 4
// NEED to subtract 2^4 -1 = 15

wire [8-1 : 0] bias;

assign bias =  ((1<< (8 -1)) -1);

	assign RoundE = NormE - 9'd15 - 9'd15 + 9'd127 ;
	assign RoundEP = NormE - 9'd15 - 9'd15 + 9'd127 ;
	assign RoundM = NormM ;
	assign RoundMP = NormM ;

endmodule

module FPMult_RoundModule_dspchain(
		RoundM,
		RoundMP,
		RoundE,
		RoundEP,
		Sp,
		GRS,
		InputExc,
		Z,
		Flags
    );

	// Input Ports
	input [23:0] RoundM ;									// Normalized 10
	input [23:0] RoundMP ;									// Normalized 5
	input [8:0] RoundE ;									// Normalized 10 + 1
	input [8:0] RoundEP ;									// Normalized 5 + 1
	input Sp ;												// Product sign
	input GRS ;
	input [4:0] InputExc ;
	
	// Output Ports
	output [32-1:0] Z ;										// Final product
	output [4:0] Flags ;
	
	// Internal Signals
	wire [8:0] FinalE ;									// Rounded 5
	wire [23:0] FinalM;
	wire [23:0] PreShiftM;
	
	assign PreShiftM = GRS ? RoundMP : RoundM ;	// Round up if R and (G or S)
	
	// Post rounding normalization (potential one bit shift> use shifted 10 if there is overflow)
	assign FinalM = (PreShiftM[23] ? {1'b0, PreShiftM[23:1]} : PreShiftM[23:0]) ;
	assign FinalE = (PreShiftM[23] ? RoundEP : RoundE) ; // Increment 5 if a shift was done
	
	
	assign Z = {Sp, FinalE[8-1:0], FinalM[21-1:0], 2'b0} ;   // Putting the pieces together
	assign Flags = InputExc[4:0];

endmodule


module FPAddSub_single_dspchain(
		clk,
		rst,
		a,
		b,
		operation,
		result,
		flags
	);

// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [31:0] a ;								// Input A, a 32-bit floating point number
	input [31:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [31:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754

	reg [68:0]pipe_1;
	reg [54:0]pipe_2;
	reg [45:0]pipe_3;


//internal module wires

//output ports
	wire Opout;
	wire Sa;
	wire Sb;
	wire MaxAB;
	wire [7:0] CExp;
	wire [4:0] Shift;
	wire [22:0] Mmax;
	wire [4:0] InputExc;
	wire [23:0] Mmin_3;

	wire [32:0] SumS_5 ;
	wire [4:0] Shift_1;							
	wire PSgn ;							
	wire Opr ;	
	
	wire [22:0] NormM ;				// Normalized mantissa
	wire [8:0] NormE ;					// Adjusted exponent
	wire ZeroSum ;						// Zero flag
	wire NegE ;							// Flag indicating negative exponent
	wire R ;								// Round bit
	wire S ;								// Final sticky bit
	wire FG ;

FPAddSub_a_dspchain M1(a,b,operation,Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3);

FpAddSub_b_dspchain M2(pipe_1[51:29],pipe_1[23:0],pipe_1[67],pipe_1[66],pipe_1[65],pipe_1[68],SumS_5,Shift_1,PSgn,Opr);

FPAddSub_c_dspchain M3(pipe_2[54:22],pipe_2[21:17],pipe_2[16:9],NormM,NormE,ZeroSum,NegE,R,S,FG);

FPAddSub_d_dspchain M4(pipe_3[13],pipe_3[22:14],pipe_3[45:23],pipe_3[11],pipe_3[10],pipe_3[9],pipe_3[8],pipe_3[7],pipe_3[6],pipe_3[5],pipe_3[12],pipe_3[4:0],result,flags );


always @ (posedge clk) begin	
		if(rst) begin
			pipe_1 <= 0;
			pipe_2 <= 0;
			pipe_3 <= 0;
		end 
		else begin
/*
pipe_1:
	[68] Opout;
	[67] Sa;
	[66] Sb;
	[65] MaxAB;
	[64:57] CExp;
	[56:52] Shift;
	[51:29] Mmax;
	[28:24] InputExc;
	[23:0] Mmin_3;	
*/

pipe_1 <= {Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3};

/*
pipe_2:
	[54:22]SumS_5;
	[21:17]Shift;
	[16:9]CExp;	
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_2 <= {SumS_5,Shift_1,pipe_1[64:57], pipe_1[67], pipe_1[66], pipe_1[68], pipe_1[65], pipe_1[28:24] };

/*
pipe_3:
	[45:23] NormM ;				
	[22:14] NormE ;					
	[13]ZeroSum ;						
	[12]NegE ;							
	[11]R ;								
	[10]S ;								
	[9]FG ;
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_3 <= {NormM,NormE,ZeroSum,NegE,R,S,FG, pipe_2[8], pipe_2[7], pipe_2[6], pipe_2[5], pipe_2[4:0] };

end
end

endmodule

// Prealign + Align + Shift 1 + Shift 2
module FPAddSub_a_dspchain(
		A,
		B,
		operation,
		Opout,
		Sa,
		Sb,
		MaxAB,
		CExp,
		Shift,
		Mmax,
		InputExc,
		Mmin_3
		
		
	);
	
	// Input ports
	input [31:0] A ;										// Input A, a 32-bit floating point number
	input [31:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	//output ports
	output Opout;
	output Sa;
	output Sb;
	output MaxAB;
	output [7:0] CExp;
	output [4:0] Shift;
	output [22:0] Mmax;
	output [4:0] InputExc;
	output [23:0] Mmin_3;	
							
	wire [9:0] ShiftDet ;							
	wire [30:0] Aout ;
	wire [30:0] Bout ;
	

	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [7:0] DAB ;										// ExpA - ExpB					
	wire [7:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[30:23]) & |(A[22:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[30:23]) & |(B[22:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[30:23]) & ~|(A[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[30:23]) & ~|(B[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
  assign DAB = (A[30:23] + ~(B[30:23]) + 1) ;
	assign DBA = (B[30:23] + ~(A[30:23]) + 1) ;

	assign Sa = A[31] ;									// A's sign bit
	assign Sb = B[31] ;									// B's sign	bit
	assign ShiftDet = {DBA[4:0], DAB[4:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[30:0] ;
	assign Bout = B[30:0] ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Output ports
													// Number of steps to smaller mantissa shift right
	wire [22:0] Mmin_1 ;							// Smaller mantissa 
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (Aout[30:0] < Bout[30:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[9:5] : ShiftDet[4:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin_1 = MaxAB ? Aout[22:0] : Bout[22:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? Bout[22:0]: Aout[22:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? Bout[30:23] : Aout[30:23]) ;	

// Input ports
					// Smaller mantissa after 16|12|8|4 shift
	wire [2:0] Shift_1 ;						// Shift amount
	
	assign Shift_1 = Shift [4:2];

	wire [23:0] Mmin_2 ;						// The smaller mantissa
	
	// Internal signals
	reg	  [23:0]		Lvl1;
	reg	  [23:0]		Lvl2;
	wire    [47:0]    Stage1;	
	integer           i;                // Loop variable
	
	always @(*) begin						
		// Rotate by 16?
		Lvl1 <= Shift_1[2] ? {17'b00000000000000001, Mmin_1[22:16]} : {1'b1, Mmin_1}; 
	end
	
	assign Stage1 = {Lvl1, Lvl1};
	
	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift_1[1:0])
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[23:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[23:19] <= 0; end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end Lvl2[23:15] <= 0; end
			// Rotate by 12	
			2'b11:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[23:11] <= 0; end
	  endcase
	end
	
	// Assign output to next shift stage
	assign Mmin_2 = Lvl2;
								// Smaller mantissa after 16|12|8|4 shift
	wire [1:0] Shift_2 ;						// Shift amount
	
	assign Shift_2 =Shift  [1:0] ;
					// The smaller mantissa
	
	// Internal Signal
	reg	  [23:0]		Lvl3;
	wire    [47:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {Mmin_2, Mmin_2};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_2[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[23:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end Lvl3[23] <= 0; end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end Lvl3[23:22] <= 0; end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end Lvl3[23:21] <= 0; end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin_3 = Lvl3;	

	
endmodule

module FpAddSub_b_dspchain(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		SumS_5,
		Shift,
		PSgn,
		Opr
);
	input [22:0] Mmax ;					// The larger mantissa
	input [23:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	wire [32:0] Sum ;	
						// Output ports
	output [32:0] SumS_5 ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount				// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation

	// Perform effective operation
	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, 8'b00000000} - {Mmin, 8'b00000000}) : ({1'b1, Mmax, 8'b00000000} + {Mmin, 8'b00000000}) ;
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

		// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[32] ? 5'b00000 :	 
		Sum[31] ? 5'b00001 : 
		Sum[30] ? 5'b00010 : 
		Sum[29] ? 5'b00011 : 
		Sum[28] ? 5'b00100 : 
		Sum[27] ? 5'b00101 : 
		Sum[26] ? 5'b00110 : 
		Sum[25] ? 5'b00111 :
		Sum[24] ? 5'b01000 :
		Sum[23] ? 5'b01001 :
		Sum[22] ? 5'b01010 :
		Sum[21] ? 5'b01011 :
		Sum[20] ? 5'b01100 :
		Sum[19] ? 5'b01101 :
		Sum[18] ? 5'b01110 :
		Sum[17] ? 5'b01111 :
		Sum[16] ? 5'b10000 :
		Sum[15] ? 5'b10001 :
		Sum[14] ? 5'b10010 :
		Sum[13] ? 5'b10011 :
		Sum[12] ? 5'b10100 :
		Sum[11] ? 5'b10101 :
		Sum[10] ? 5'b10110 :
		Sum[9] ? 5'b10111 :
		Sum[8] ? 5'b11000 :
		Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [32:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[16:0], 16'b0000000000000000} : Sum; 
	end
	
	// Assign outputs
	assign SumS_5 = Lvl1;	

endmodule

module FPAddSub_c_dspchain(
		SumS_5,
		Shift,
		CExp,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [32:0] SumS_5 ;						// Smaller mantissa after 16|12|8|4 shift
	
	input [4:0] Shift ;						// Shift amount
	
// Input ports
	
	input [7:0] CExp ;
	

	// Output ports
	output [22:0] NormM ;				// Normalized mantissa
	output [8:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;


	wire [3:0]Shift_1;
	assign Shift_1 = Shift [3:0];
	// Output ports
	wire [32:0] SumS_7 ;						// The smaller mantissa
	
	reg	  [32:0]		Lvl2;
	wire    [65:0]    Stage1;	
	reg	  [32:0]		Lvl3;
	wire    [65:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {SumS_5, SumS_5};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: Lvl2 <= Stage1[32:0];       		
			// Rotate by 4
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
			// Rotate by 8
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
			// Rotate by 12
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_1[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[32:0];
			// Rotate by 1
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
			// Rotate by 2
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
			// Rotate by 3
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
	  endcase
	end
	
	// Assign outputs
	assign SumS_7 = Lvl3;						// Take out smaller mantissa



	
	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [8:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [8:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = SumS_7[32] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|SumS_7 ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[8] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = SumS_7[31:9] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = SumS_7[8] ; 
	assign R = SumS_7[7] ;
	assign S = |SumS_7[6:0] ;		
	
endmodule

module FPAddSub_d_dspchain(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		NegE,
		InputExc,
		P,
		Flags 
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [8:0] NormE ;				// Normalized exponent
	input [22:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	

	input NegE ;						// Negative exponent?
	input [4:0] InputExc ;					// Exceptions in inputs A and B

	// Output ports
	output [31:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// 
	wire [31:0] Z ;					// Final result
	wire EOF ;
	
	// Internal signals
	wire [23:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [22:0] RoundM ;				// The final rounded sum
	wire [8:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	wire FSgn;
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[22:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[23] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? 8'b00000000 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[7:0], RoundM[22:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[8];

/////////////////////////////////////////////////////////////////////////////////////////////////////////



	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[30:23]) & ~|(Z[30:23]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule

`endif 


module dbram_2048_40bit (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b,reset
); 

parameter AWIDTH=11;
parameter NUM_WORDS=2048;
parameter DWIDTH=40;
input clk, reset;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

reg count; 

always@(posedge clk) begin 

if (reset) begin 
	count <= 1'b0; 
end
else begin 
	count <= ~count; 
end

end

wire [(AWIDTH-1):0] address_a1,address_a2;
wire [(AWIDTH-1):0] address_b1,address_b2;
wire  wren_a1,wren_a2;
wire  wren_b1,wren_b2;
wire [(DWIDTH-1):0] data_a1,data_a2;
wire [(DWIDTH-1):0] data_b1,data_b2;
wire [(DWIDTH-1):0] out_a1,out_a2;
wire [(DWIDTH-1):0] out_b1,out_b2;

assign address_a1 = count|address_a; 
assign address_a2 = (~count)|address_a;
assign address_b1 = count|address_b; 
assign address_b2 = (~count)|address_b;
assign wren_a1 = count|wren_a; 
assign wren_a2 = (~count)|wren_a; 
assign wren_b1 = count|wren_b; 
assign wren_b2 = (~count)|wren_b; 
assign data_a1 = count|data_a;
assign data_a2 = (~count)|data_a;
assign data_b1 = count|data_b;
assign data_b2 = (~count)|data_b;
always@(posedge clk) begin 
out_a <= count?out_a1:out_a2;
out_b <= count?out_b1:out_b2;
end
dpram_2048_40bit_db inst1(.clk(clk),.address_a(address_a1),.address_b(address_b1),.wren_a(wren_a1),.wren_b(wren_b1),.data_a(data_a1),.data_b(data_b1),.out_a(out_a1),.out_b(out_b1));
dpram_2048_40bit_db inst2(.clk(clk),.address_a(address_a2),.address_b(address_b2),.wren_a(wren_a2),.wren_b(wren_b2),.data_a(data_a2),.data_b(data_b2),.out_a(out_a2),.out_b(out_b2));


endmodule

module dpram_2048_40bit_db (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b
);
parameter AWIDTH=11;
parameter NUM_WORDS=2048;
parameter DWIDTH=40;
input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren_a) 
      ram[address_a] <= data_a;
  if (wren_b) 
      ram[address_b] <= data_b;
  out_a <= ram[address_a];
  out_b <= ram[address_b];
end
  

`else

defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

dual_port_ram u_dual_port_ram(
.addr1(address_a),
.we1(wren_a),
.data1(data_a),
.out1(out_a),
.addr2(address_b),
.we2(wren_b),
.data2(data_b),
.out2(out_b),
.clk(clk)
);

`endif
endmodule

`timescale 1ns / 1ps
//`define complex_dsp
`define DWIDTH 16
`define AWIDTH 10
`define MEM_SIZE 1024

`define MAT_MUL_SIZE 4
`define MASK_WIDTH 4
`define LOG2_MAT_MUL_SIZE 2

`define NUM_CYCLES_IN_MAC 3
`define MEM_ACCESS_LATENCY 1
`define REG_DATAWIDTH 32
`define REG_ADDRWIDTH 8
`define ADDR_STRIDE_WIDTH 10
`define MAX_BITS_POOL 3
`define EXPONENT 5
`define MANTISSA 10
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/10/2020 11:43:24 PM
// Design Name: 
// Module Name: matmul_4x4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module matmul_4x4_fp_systolic(
 clk,
 reset,
 pe_reset,
 start_mat_mul,
 done_mat_mul,
 address_mat_a,
 address_mat_b,
 address_mat_c,
 address_stride_a,
 address_stride_b,
 address_stride_c,
 a_data,
 b_data,
 a_data_in, //Data values coming in from previous matmul - systolic connections
 b_data_in,
 c_data_in, //Data values coming in from previous matmul - systolic shifting
 c_data_out, //Data values going out to next matmul - systolic shifting
 a_data_out,
 b_data_out,
 a_addr,
 b_addr,
 c_addr,
 c_data_available,
 validity_mask_a_rows,
 validity_mask_a_cols_b_rows,
 validity_mask_b_cols,
 final_mat_mul_size,
 a_loc,
 b_loc
);

 input clk;
 input reset;
 input pe_reset;
 input start_mat_mul;
 output done_mat_mul;
 input [`AWIDTH-1:0] address_mat_a;
 input [`AWIDTH-1:0] address_mat_b;
 input [`AWIDTH-1:0] address_mat_c;
 input [`ADDR_STRIDE_WIDTH-1:0] address_stride_a;
 input [`ADDR_STRIDE_WIDTH-1:0] address_stride_b;
 input [`ADDR_STRIDE_WIDTH-1:0] address_stride_c;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_in;
 output [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out;
 output [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data_out;
 output [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data_out;
 output [`AWIDTH-1:0] a_addr;
 output [`AWIDTH-1:0] b_addr;
 output [`AWIDTH-1:0] c_addr;
 output c_data_available;
 input [`MASK_WIDTH-1:0] validity_mask_a_rows;
 input [`MASK_WIDTH-1:0] validity_mask_a_cols_b_rows;
 input [`MASK_WIDTH-1:0] validity_mask_b_cols;
//7:0 is okay here. We aren't going to make a matmul larger than 128x128
//In fact, these will get optimized out by the synthesis tool, because
//we hardcode them at the instantiation level.
 input [7:0] final_mat_mul_size;
 input [7:0] a_loc;
 input [7:0] b_loc;

//////////////////////////////////////////////////////////////////////////
// Logic for clock counting and when to assert done
//////////////////////////////////////////////////////////////////////////

reg done_mat_mul;
//This is 7 bits because the expectation is that clock count will be pretty
//small. For large matmuls, this will need to increased to have more bits.
//In general, a systolic multiplier takes 4*N-2+P cycles, where N is the size 
//of the matmul and P is the number of pipleine stages in the MAC block.
reg [7:0] clk_cnt;

//Finding out number of cycles to assert matmul done.
//When we have to save the outputs to accumulators, then we don't need to
//shift out data. So, we can assert done_mat_mul early.
//In the normal case, we have to include the time to shift out the results. 
//Note: the count expression used to contain "4*final_mat_mul_size", but 
//to avoid multiplication, we now use "final_mat_mul_size<<2"
wire [7:0] clk_cnt_for_done;
assign clk_cnt_for_done = 
                          ((final_mat_mul_size<<2) - 2 + `NUM_CYCLES_IN_MAC) ;  

always @(posedge clk) begin
  if (reset || ~start_mat_mul) begin
    clk_cnt <= 0;
    done_mat_mul <= 0;
  end
  else if (clk_cnt == clk_cnt_for_done) begin
    done_mat_mul <= 1;
    clk_cnt <= clk_cnt + 1;
  end
  else if (done_mat_mul == 0) begin
    clk_cnt <= clk_cnt + 1;
  end    
  else begin
    done_mat_mul <= 0;
    clk_cnt <= clk_cnt + 1;
  end
end


wire [`DWIDTH-1:0] a0_data;
wire [`DWIDTH-1:0] a1_data;
wire [`DWIDTH-1:0] a2_data;
wire [`DWIDTH-1:0] a3_data;
wire [`DWIDTH-1:0] b0_data;
wire [`DWIDTH-1:0] b1_data;
wire [`DWIDTH-1:0] b2_data;
wire [`DWIDTH-1:0] b3_data;
wire [`DWIDTH-1:0] a1_data_delayed_1;
wire [`DWIDTH-1:0] a2_data_delayed_1;
wire [`DWIDTH-1:0] a2_data_delayed_2;
wire [`DWIDTH-1:0] a3_data_delayed_1;
wire [`DWIDTH-1:0] a3_data_delayed_2;
wire [`DWIDTH-1:0] a3_data_delayed_3;
wire [`DWIDTH-1:0] b1_data_delayed_1;
wire [`DWIDTH-1:0] b2_data_delayed_1;
wire [`DWIDTH-1:0] b2_data_delayed_2;
wire [`DWIDTH-1:0] b3_data_delayed_1;
wire [`DWIDTH-1:0] b3_data_delayed_2;
wire [`DWIDTH-1:0] b3_data_delayed_3;

//////////////////////////////////////////////////////////////////////////
// Instantiation of systolic data setup
//////////////////////////////////////////////////////////////////////////
systolic_data_setup_systolic_4x4_fp u_systolic_data_setup_systolic_4x4_fp(
.clk(clk),
.reset(reset),
.start_mat_mul(start_mat_mul),
.a_addr(a_addr),
.b_addr(b_addr),
.address_mat_a(address_mat_a),
.address_mat_b(address_mat_b),
.address_stride_a(address_stride_a),
.address_stride_b(address_stride_b),
.a_data(a_data),
.b_data(b_data),
.clk_cnt(clk_cnt),
.a0_data(a0_data),
.a1_data_delayed_1(a1_data_delayed_1),
.a2_data_delayed_2(a2_data_delayed_2),
.a3_data_delayed_3(a3_data_delayed_3),
.b0_data(b0_data),
.b1_data_delayed_1(b1_data_delayed_1),
.b2_data_delayed_2(b2_data_delayed_2),
.b3_data_delayed_3(b3_data_delayed_3),
.validity_mask_a_rows(validity_mask_a_rows),
.validity_mask_a_cols_b_rows(validity_mask_a_cols_b_rows),
.validity_mask_b_cols(validity_mask_b_cols),
.final_mat_mul_size(final_mat_mul_size),
.a_loc(a_loc),
.b_loc(b_loc)
);


//////////////////////////////////////////////////////////////////////////
// Logic to mux data_in coming from neighboring matmuls
//////////////////////////////////////////////////////////////////////////
wire [`DWIDTH-1:0] a0;
wire [`DWIDTH-1:0] a1;
wire [`DWIDTH-1:0] a2;
wire [`DWIDTH-1:0] a3;
wire [`DWIDTH-1:0] b0;
wire [`DWIDTH-1:0] b1;
wire [`DWIDTH-1:0] b2;
wire [`DWIDTH-1:0] b3;

wire [`DWIDTH-1:0] a0_data_in;
wire [`DWIDTH-1:0] a1_data_in;
wire [`DWIDTH-1:0] a2_data_in;
wire [`DWIDTH-1:0] a3_data_in;
assign a0_data_in = a_data_in[`DWIDTH-1:0];
assign a1_data_in = a_data_in[2*`DWIDTH-1:`DWIDTH];
assign a2_data_in = a_data_in[3*`DWIDTH-1:2*`DWIDTH];
assign a3_data_in = a_data_in[4*`DWIDTH-1:3*`DWIDTH];

wire [`DWIDTH-1:0] b0_data_in;
wire [`DWIDTH-1:0] b1_data_in;
wire [`DWIDTH-1:0] b2_data_in;
wire [`DWIDTH-1:0] b3_data_in;
assign b0_data_in = b_data_in[`DWIDTH-1:0];
assign b1_data_in = b_data_in[2*`DWIDTH-1:`DWIDTH];
assign b2_data_in = b_data_in[3*`DWIDTH-1:2*`DWIDTH];
assign b3_data_in = b_data_in[4*`DWIDTH-1:3*`DWIDTH];

//If b_loc is 0, that means this matmul block is on the top-row of the
//final large matmul. In that case, b will take inputs from mem.
//If b_loc != 0, that means this matmul block is not on the top-row of the
//final large matmul. In that case, b will take inputs from the matmul on top
//of this one.
assign a0 = (b_loc==0) ? a0_data           : a0_data_in;
assign a1 = (b_loc==0) ? a1_data_delayed_1 : a1_data_in;
assign a2 = (b_loc==0) ? a2_data_delayed_2 : a2_data_in;
assign a3 = (b_loc==0) ? a3_data_delayed_3 : a3_data_in;

//If a_loc is 0, that means this matmul block is on the left-col of the
//final large matmul. In that case, a will take inputs from mem.
//If a_loc != 0, that means this matmul block is not on the left-col of the
//final large matmul. In that case, a will take inputs from the matmul on left
//of this one.
assign b0 = (a_loc==0) ? b0_data           : b0_data_in;
assign b1 = (a_loc==0) ? b1_data_delayed_1 : b1_data_in;
assign b2 = (a_loc==0) ? b2_data_delayed_2 : b2_data_in;
assign b3 = (a_loc==0) ? b3_data_delayed_3 : b3_data_in;


wire [`DWIDTH-1:0] matrixC00;
wire [`DWIDTH-1:0] matrixC01;
wire [`DWIDTH-1:0] matrixC02;
wire [`DWIDTH-1:0] matrixC03;
wire [`DWIDTH-1:0] matrixC10;
wire [`DWIDTH-1:0] matrixC11;
wire [`DWIDTH-1:0] matrixC12;
wire [`DWIDTH-1:0] matrixC13;
wire [`DWIDTH-1:0] matrixC20;
wire [`DWIDTH-1:0] matrixC21;
wire [`DWIDTH-1:0] matrixC22;
wire [`DWIDTH-1:0] matrixC23;
wire [`DWIDTH-1:0] matrixC30;
wire [`DWIDTH-1:0] matrixC31;
wire [`DWIDTH-1:0] matrixC32;
wire [`DWIDTH-1:0] matrixC33;


//////////////////////////////////////////////////////////////////////////
// Instantiation of the output logic
//////////////////////////////////////////////////////////////////////////
output_logic_systolic_4x4_fp u_output_logic_systolic_4x4_fp(
.clk(clk),
.reset(reset),
.start_mat_mul(start_mat_mul),
.done_mat_mul(done_mat_mul),
.address_mat_c(address_mat_c),
.address_stride_c(address_stride_c),
.c_data_out(c_data_out),
.c_data_in(c_data_in),
.c_addr(c_addr),
.c_data_available(c_data_available),
.clk_cnt(clk_cnt),
.final_mat_mul_size(final_mat_mul_size),
.matrixC00(matrixC00),
.matrixC01(matrixC01),
.matrixC02(matrixC02),
.matrixC03(matrixC03),
.matrixC10(matrixC10),
.matrixC11(matrixC11),
.matrixC12(matrixC12),
.matrixC13(matrixC13),
.matrixC20(matrixC20),
.matrixC21(matrixC21),
.matrixC22(matrixC22),
.matrixC23(matrixC23),
.matrixC30(matrixC30),
.matrixC31(matrixC31),
.matrixC32(matrixC32),
.matrixC33(matrixC33)
);

//////////////////////////////////////////////////////////////////////////
// Instantiations of the actual PEs
//////////////////////////////////////////////////////////////////////////
systolic_pe_matrix_systolic_4x4_fp u_systolic_pe_matrix_systolic_4x4_fp(
.reset(reset),
.clk(clk),
.pe_reset(pe_reset),
.start_mat_mul(start_mat_mul),
.a0(a0), 
.a1(a1), 
.a2(a2), 
.a3(a3),
.b0(b0), 
.b1(b1), 
.b2(b2), 
.b3(b3),
.matrixC00(matrixC00),
.matrixC01(matrixC01),
.matrixC02(matrixC02),
.matrixC03(matrixC03),
.matrixC10(matrixC10),
.matrixC11(matrixC11),
.matrixC12(matrixC12),
.matrixC13(matrixC13),
.matrixC20(matrixC20),
.matrixC21(matrixC21),
.matrixC22(matrixC22),
.matrixC23(matrixC23),
.matrixC30(matrixC30),
.matrixC31(matrixC31),
.matrixC32(matrixC32),
.matrixC33(matrixC33),
.a_data_out(a_data_out),
.b_data_out(b_data_out)
);

endmodule

//////////////////////////////////////////////////////////////////////////
// Output logic
//////////////////////////////////////////////////////////////////////////
module output_logic_systolic_4x4_fp(
clk,
reset,
start_mat_mul,
done_mat_mul,
address_mat_c,
address_stride_c,
c_data_in,
c_data_out, //Data values going out to next matmul - systolic shifting
c_addr,
c_data_available,
clk_cnt,
final_mat_mul_size,
matrixC00,
matrixC01,
matrixC02,
matrixC03,
matrixC10,
matrixC11,
matrixC12,
matrixC13,
matrixC20,
matrixC21,
matrixC22,
matrixC23,
matrixC30,
matrixC31,
matrixC32,
matrixC33
);

input clk;
input reset;
input start_mat_mul;
input done_mat_mul;
input [`AWIDTH-1:0] address_mat_c;
input [`ADDR_STRIDE_WIDTH-1:0] address_stride_c;
input [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_in;
output [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out;
output [`AWIDTH-1:0] c_addr;
output c_data_available;
input [7:0] clk_cnt;
//output row_latch_en;
input [7:0] final_mat_mul_size;
input [`DWIDTH-1:0] matrixC00;
input [`DWIDTH-1:0] matrixC01;
input [`DWIDTH-1:0] matrixC02;
input [`DWIDTH-1:0] matrixC03;
input [`DWIDTH-1:0] matrixC10;
input [`DWIDTH-1:0] matrixC11;
input [`DWIDTH-1:0] matrixC12;
input [`DWIDTH-1:0] matrixC13;
input [`DWIDTH-1:0] matrixC20;
input [`DWIDTH-1:0] matrixC21;
input [`DWIDTH-1:0] matrixC22;
input [`DWIDTH-1:0] matrixC23;
input [`DWIDTH-1:0] matrixC30;
input [`DWIDTH-1:0] matrixC31;
input [`DWIDTH-1:0] matrixC32;
input [`DWIDTH-1:0] matrixC33;

wire row_latch_en;

//////////////////////////////////////////////////////////////////////////
// Logic to capture matrix C data from the PEs and shift it out
//////////////////////////////////////////////////////////////////////////

//assign row_latch_en = (clk_cnt==(`MAT_MUL_SIZE + (a_loc+b_loc) * `BB_MAT_MUL_SIZE + 10 +  `NUM_CYCLES_IN_MAC - 1));
//Writing the line above to avoid multiplication:
//assign row_latch_en = (clk_cnt==(`MAT_MUL_SIZE + ((a_loc+b_loc) << `LOG2_MAT_MUL_SIZE) + 10 +  `NUM_CYCLES_IN_MAC - 1));
//Fixing bug. The line above is inaccurate. Using the line below. 
//TODO: This line needs to be fixed to include a_loc and b_loc ie. when final_mat_mul_size is different from `MAT_MUL_SIZE
assign row_latch_en =  
                       //((clk_cnt == ((`MAT_MUL_SIZE<<2) - `MAT_MUL_SIZE -2 +`NUM_CYCLES_IN_MAC)));
                       ((clk_cnt == ((final_mat_mul_size<<2) - final_mat_mul_size -1 +`NUM_CYCLES_IN_MAC)));

reg c_data_available;
reg [`AWIDTH-1:0] c_addr;
reg start_capturing_c_data;
integer counter;
reg [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out;
reg [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out_1;
reg [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out_2;
reg [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out_3;

wire [`MAT_MUL_SIZE*`DWIDTH-1:0] col0;
wire [`MAT_MUL_SIZE*`DWIDTH-1:0] col1;
wire [`MAT_MUL_SIZE*`DWIDTH-1:0] col2;
wire [`MAT_MUL_SIZE*`DWIDTH-1:0] col3;
assign col0 = {matrixC30, matrixC20, matrixC10, matrixC00};
assign col1 = {matrixC31, matrixC21, matrixC11, matrixC01};
assign col2 = {matrixC32, matrixC22, matrixC12, matrixC02};
assign col3 = {matrixC33, matrixC23, matrixC13, matrixC03};

//If save_output_to_accum is asserted, that means we are not intending to shift
//out the outputs, because the outputs are still partial sums. 
wire condition_to_start_shifting_output;
assign condition_to_start_shifting_output = 
                          row_latch_en ;  

//For larger matmuls, this logic will have more entries in the case statement
always @(posedge clk) begin
  if (reset | ~start_mat_mul) begin
    start_capturing_c_data <= 1'b0;
    c_data_available <= 1'b0;
    c_addr <= address_mat_c+address_stride_c;
    c_data_out <= 0;
    counter <= 0;
    c_data_out_1 <= 0; 
    c_data_out_2 <= 0; 
    c_data_out_3 <= 0; 
  end
  else if (condition_to_start_shifting_output) begin
    start_capturing_c_data <= 1'b1;
    c_data_available <= 1'b1;
    c_addr <= c_addr - address_stride_c;
    c_data_out <= col0; 
    c_data_out_1 <= col1; 
    c_data_out_2 <= col2; 
    c_data_out_3 <= col3; 
    counter <= counter + 1;
  end 
  else if (done_mat_mul) begin
    start_capturing_c_data <= 1'b0;
    c_data_available <= 1'b0;
    c_addr <= address_mat_c+address_stride_c;
    c_data_out <= 0;
    c_data_out_1 <= 0;
    c_data_out_2 <= 0;
    c_data_out_3 <= 0;
  end 
  else if (counter >= `MAT_MUL_SIZE) begin
    c_addr <= c_addr - address_stride_c;
    c_data_out <= c_data_out_1;
    c_data_out_1 <= c_data_out_2;
    c_data_out_2 <= c_data_out_3;
    c_data_out_3 <= c_data_in;
  end
  else if (start_capturing_c_data) begin
    c_data_available <= 1'b1;
    c_addr <= c_addr - address_stride_c;
    counter <= counter + 1;
    c_data_out <= c_data_out_1;
    c_data_out_1 <= c_data_out_2;
    c_data_out_2 <= c_data_out_3;
    c_data_out_3 <= c_data_in;
  end
end

endmodule

//////////////////////////////////////////////////////////////////////////
// Systolic data setup
//////////////////////////////////////////////////////////////////////////
module systolic_data_setup_systolic_4x4_fp(
clk,
reset,
start_mat_mul,
a_addr,
b_addr,
address_mat_a,
address_mat_b,
address_stride_a,
address_stride_b,
a_data,
b_data,
clk_cnt,
a0_data,
a1_data_delayed_1,
a2_data_delayed_2,
a3_data_delayed_3,
b0_data,
b1_data_delayed_1,
b2_data_delayed_2,
b3_data_delayed_3,
validity_mask_a_rows,
validity_mask_a_cols_b_rows,
validity_mask_b_cols,
final_mat_mul_size,
a_loc,
b_loc
);

input clk;
input reset;
input start_mat_mul;
output [`AWIDTH-1:0] a_addr;
output [`AWIDTH-1:0] b_addr;
input [`AWIDTH-1:0] address_mat_a;
input [`AWIDTH-1:0] address_mat_b;
input [`ADDR_STRIDE_WIDTH-1:0] address_stride_a;
input [`ADDR_STRIDE_WIDTH-1:0] address_stride_b;
input [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data;
input [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data;
input [7:0] clk_cnt;
output [`DWIDTH-1:0] a0_data;
output [`DWIDTH-1:0] a1_data_delayed_1;
output [`DWIDTH-1:0] a2_data_delayed_2;
output [`DWIDTH-1:0] a3_data_delayed_3;
output [`DWIDTH-1:0] b0_data;
output [`DWIDTH-1:0] b1_data_delayed_1;
output [`DWIDTH-1:0] b2_data_delayed_2;
output [`DWIDTH-1:0] b3_data_delayed_3;
input [`MASK_WIDTH-1:0] validity_mask_a_rows;
input [`MASK_WIDTH-1:0] validity_mask_a_cols_b_rows;
input [`MASK_WIDTH-1:0] validity_mask_b_cols;
input [7:0] final_mat_mul_size;
input [7:0] a_loc;
input [7:0] b_loc;

wire [`DWIDTH-1:0] a0_data;
wire [`DWIDTH-1:0] a1_data;
wire [`DWIDTH-1:0] a2_data;
wire [`DWIDTH-1:0] a3_data;
wire [`DWIDTH-1:0] b0_data;
wire [`DWIDTH-1:0] b1_data;
wire [`DWIDTH-1:0] b2_data;
wire [`DWIDTH-1:0] b3_data;

//////////////////////////////////////////////////////////////////////////
// Logic to generate addresses to BRAM A
//////////////////////////////////////////////////////////////////////////
reg [`AWIDTH-1:0] a_addr;
reg a_mem_access; //flag that tells whether the matmul is trying to access memory or not

always @(posedge clk) begin
  //else if (clk_cnt >= a_loc*`MAT_MUL_SIZE+final_mat_mul_size) begin
  //Writing the line above to avoid multiplication:
  if ((reset || ~start_mat_mul) || (clk_cnt >= (a_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
      a_addr <= address_mat_a-address_stride_a;
    a_mem_access <= 0;
  end

  //else if ((clk_cnt >= a_loc*`MAT_MUL_SIZE) && (clk_cnt < a_loc*`MAT_MUL_SIZE+final_mat_mul_size)) begin
  //Writing the line above to avoid multiplication:
  else if ((clk_cnt >= (a_loc<<`LOG2_MAT_MUL_SIZE)) && (clk_cnt < (a_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
      a_addr <= a_addr + address_stride_a;
    a_mem_access <= 1;
  end
end  

//////////////////////////////////////////////////////////////////////////
// Logic to generate valid signals for data coming from BRAM A
//////////////////////////////////////////////////////////////////////////
reg [7:0] a_mem_access_counter;
always @(posedge clk) begin
  if (reset || ~start_mat_mul) begin
    a_mem_access_counter <= 0;
  end
  else if (a_mem_access == 1) begin
    a_mem_access_counter <= a_mem_access_counter + 1;  

  end
  else begin
    a_mem_access_counter <= 0;
  end
end

wire a_data_valid; //flag that tells whether the data from memory is valid
assign a_data_valid = 
       ((validity_mask_a_cols_b_rows[0]==1'b0 && a_mem_access_counter==1) ||
        (validity_mask_a_cols_b_rows[1]==1'b0 && a_mem_access_counter==2) ||
        (validity_mask_a_cols_b_rows[2]==1'b0 && a_mem_access_counter==3) ||
        (validity_mask_a_cols_b_rows[3]==1'b0 && a_mem_access_counter==4)) ?
        1'b0 : (a_mem_access_counter >= `MEM_ACCESS_LATENCY);

//////////////////////////////////////////////////////////////////////////
// Logic to delay certain parts of the data received from BRAM A (systolic data setup)
//////////////////////////////////////////////////////////////////////////
//Slice data into chunks and qualify it with whether it is valid or not
assign a0_data = a_data[`DWIDTH-1:0] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[0]}};
assign a1_data = a_data[2*`DWIDTH-1:`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[1]}};
assign a2_data = a_data[3*`DWIDTH-1:2*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[2]}};
assign a3_data = a_data[4*`DWIDTH-1:3*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[3]}};

//For larger matmuls, more such delaying flops will be needed
reg [`DWIDTH-1:0] a1_data_delayed_1;
reg [`DWIDTH-1:0] a2_data_delayed_1;
reg [`DWIDTH-1:0] a2_data_delayed_2;
reg [`DWIDTH-1:0] a3_data_delayed_1;
reg [`DWIDTH-1:0] a3_data_delayed_2;
reg [`DWIDTH-1:0] a3_data_delayed_3;
always @(posedge clk) begin
  if (reset || ~start_mat_mul || clk_cnt==0) begin
    a1_data_delayed_1 <= 0;
    a2_data_delayed_1 <= 0;
    a2_data_delayed_2 <= 0;
    a3_data_delayed_1 <= 0;
    a3_data_delayed_2 <= 0;
    a3_data_delayed_3 <= 0;
  end
  else begin
    a1_data_delayed_1 <= a1_data;
    a2_data_delayed_1 <= a2_data;
    a2_data_delayed_2 <= a2_data_delayed_1;
    a3_data_delayed_1 <= a3_data;
    a3_data_delayed_2 <= a3_data_delayed_1;
    a3_data_delayed_3 <= a3_data_delayed_2;
  end
end

//////////////////////////////////////////////////////////////////////////
// Logic to generate addresses to BRAM B
//////////////////////////////////////////////////////////////////////////
reg [`AWIDTH-1:0] b_addr;
reg b_mem_access; //flag that tells whether the matmul is trying to access memory or not

always @(posedge clk) begin
  //else if (clk_cnt >= b_loc*`MAT_MUL_SIZE+final_mat_mul_size) begin
  //Writing the line above to avoid multiplication:
  if ((reset || ~start_mat_mul) || (clk_cnt >= (b_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
      b_addr <= address_mat_b - address_stride_b;
    b_mem_access <= 0;
  end
  //else if ((clk_cnt >= b_loc*`MAT_MUL_SIZE) && (clk_cnt < b_loc*`MAT_MUL_SIZE+final_mat_mul_size)) begin
  //Writing the line above to avoid multiplication:
  else if ((clk_cnt >= (b_loc<<`LOG2_MAT_MUL_SIZE)) && (clk_cnt < (b_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
      b_addr <= b_addr + address_stride_b;
    b_mem_access <= 1;
  end
end  

//////////////////////////////////////////////////////////////////////////
// Logic to generate valid signals for data coming from BRAM B
//////////////////////////////////////////////////////////////////////////
reg [7:0] b_mem_access_counter;
always @(posedge clk) begin
  if (reset || ~start_mat_mul) begin
    b_mem_access_counter <= 0;
  end
  else if (b_mem_access == 1) begin
    b_mem_access_counter <= b_mem_access_counter + 1;  
  end
  else begin
    b_mem_access_counter <= 0;
  end
end

wire b_data_valid; //flag that tells whether the data from memory is valid
assign b_data_valid = 
       ((validity_mask_a_cols_b_rows[0]==1'b0 && b_mem_access_counter==1) ||
        (validity_mask_a_cols_b_rows[1]==1'b0 && b_mem_access_counter==2) ||
        (validity_mask_a_cols_b_rows[2]==1'b0 && b_mem_access_counter==3) ||
        (validity_mask_a_cols_b_rows[3]==1'b0 && b_mem_access_counter==4)) ?
        1'b0 : (b_mem_access_counter >= `MEM_ACCESS_LATENCY);


//////////////////////////////////////////////////////////////////////////
// Logic to delay certain parts of the data received from BRAM B (systolic data setup)
//////////////////////////////////////////////////////////////////////////
//Slice data into chunks and qualify it with whether it is valid or not
assign b0_data = b_data[`DWIDTH-1:0] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[0]}};
assign b1_data = b_data[2*`DWIDTH-1:`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[1]}};
assign b2_data = b_data[3*`DWIDTH-1:2*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[2]}};
assign b3_data = b_data[4*`DWIDTH-1:3*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[3]}};

//For larger matmuls, more such delaying flops will be needed
reg [`DWIDTH-1:0] b1_data_delayed_1;
reg [`DWIDTH-1:0] b2_data_delayed_1;
reg [`DWIDTH-1:0] b2_data_delayed_2;
reg [`DWIDTH-1:0] b3_data_delayed_1;
reg [`DWIDTH-1:0] b3_data_delayed_2;
reg [`DWIDTH-1:0] b3_data_delayed_3;
always @(posedge clk) begin
  if (reset || ~start_mat_mul || clk_cnt==0) begin
    b1_data_delayed_1 <= 0;
    b2_data_delayed_1 <= 0;
    b2_data_delayed_2 <= 0;
    b3_data_delayed_1 <= 0;
    b3_data_delayed_2 <= 0;
    b3_data_delayed_3 <= 0;
  end
  else begin
    b1_data_delayed_1 <= b1_data;
    b2_data_delayed_1 <= b2_data;
    b2_data_delayed_2 <= b2_data_delayed_1;
    b3_data_delayed_1 <= b3_data;
    b3_data_delayed_2 <= b3_data_delayed_1;
    b3_data_delayed_3 <= b3_data_delayed_2;
  end
end


endmodule



//////////////////////////////////////////////////////////////////////////
// Systolically connected PEs
//////////////////////////////////////////////////////////////////////////
module systolic_pe_matrix_systolic_4x4_fp(
reset,
clk,
pe_reset,
start_mat_mul,
a0, a1, a2, a3,
b0, b1, b2, b3,
matrixC00,
matrixC01,
matrixC02,
matrixC03,
matrixC10,
matrixC11,
matrixC12,
matrixC13,
matrixC20,
matrixC21,
matrixC22,
matrixC23,
matrixC30,
matrixC31,
matrixC32,
matrixC33,
a_data_out,
b_data_out
);

input clk;
input reset;
input pe_reset;
input start_mat_mul;
input [`DWIDTH-1:0] a0;
input [`DWIDTH-1:0] a1;
input [`DWIDTH-1:0] a2;
input [`DWIDTH-1:0] a3;
input [`DWIDTH-1:0] b0;
input [`DWIDTH-1:0] b1;
input [`DWIDTH-1:0] b2;
input [`DWIDTH-1:0] b3;
output [`DWIDTH-1:0] matrixC00;
output [`DWIDTH-1:0] matrixC01;
output [`DWIDTH-1:0] matrixC02;
output [`DWIDTH-1:0] matrixC03;
output [`DWIDTH-1:0] matrixC10;
output [`DWIDTH-1:0] matrixC11;
output [`DWIDTH-1:0] matrixC12;
output [`DWIDTH-1:0] matrixC13;
output [`DWIDTH-1:0] matrixC20;
output [`DWIDTH-1:0] matrixC21;
output [`DWIDTH-1:0] matrixC22;
output [`DWIDTH-1:0] matrixC23;
output [`DWIDTH-1:0] matrixC30;
output [`DWIDTH-1:0] matrixC31;
output [`DWIDTH-1:0] matrixC32;
output [`DWIDTH-1:0] matrixC33;
output [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data_out;
output [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data_out;

wire [`DWIDTH-1:0] a00to01, a01to02, a02to03, a03to04;
wire [`DWIDTH-1:0] a10to11, a11to12, a12to13, a13to14;
wire [`DWIDTH-1:0] a20to21, a21to22, a22to23, a23to24;
wire [`DWIDTH-1:0] a30to31, a31to32, a32to33, a33to34;

wire [`DWIDTH-1:0] b00to10, b10to20, b20to30, b30to40; 
wire [`DWIDTH-1:0] b01to11, b11to21, b21to31, b31to41;
wire [`DWIDTH-1:0] b02to12, b12to22, b22to32, b32to42;
wire [`DWIDTH-1:0] b03to13, b13to23, b23to33, b33to43;

wire effective_rst;
assign effective_rst = reset | pe_reset;

 processing_element_systolic_4x4_fp pe00(.reset(effective_rst), .clk(clk),  .in_a(a0),      .in_b(b0),  .out_a(a00to01), .out_b(b00to10), .out_c(matrixC00));
 processing_element_systolic_4x4_fp pe01(.reset(effective_rst), .clk(clk),  .in_a(a00to01), .in_b(b1),  .out_a(a01to02), .out_b(b01to11), .out_c(matrixC01));
 processing_element_systolic_4x4_fp pe02(.reset(effective_rst), .clk(clk),  .in_a(a01to02), .in_b(b2),  .out_a(a02to03), .out_b(b02to12), .out_c(matrixC02));
 processing_element_systolic_4x4_fp pe03(.reset(effective_rst), .clk(clk),  .in_a(a02to03), .in_b(b3),  .out_a(a03to04), .out_b(b03to13), .out_c(matrixC03));

 processing_element_systolic_4x4_fp pe10(.reset(effective_rst), .clk(clk),  .in_a(a1),      .in_b(b00to10), .out_a(a10to11), .out_b(b10to20), .out_c(matrixC10));
 processing_element_systolic_4x4_fp pe11(.reset(effective_rst), .clk(clk),  .in_a(a10to11), .in_b(b01to11), .out_a(a11to12), .out_b(b11to21), .out_c(matrixC11));
 processing_element_systolic_4x4_fp pe12(.reset(effective_rst), .clk(clk),  .in_a(a11to12), .in_b(b02to12), .out_a(a12to13), .out_b(b12to22), .out_c(matrixC12));
 processing_element_systolic_4x4_fp pe13(.reset(effective_rst), .clk(clk),  .in_a(a12to13), .in_b(b03to13), .out_a(a13to14), .out_b(b13to23), .out_c(matrixC13));

 processing_element_systolic_4x4_fp pe20(.reset(effective_rst), .clk(clk),  .in_a(a2),      .in_b(b10to20), .out_a(a20to21), .out_b(b20to30), .out_c(matrixC20));
 processing_element_systolic_4x4_fp pe21(.reset(effective_rst), .clk(clk),  .in_a(a20to21), .in_b(b11to21), .out_a(a21to22), .out_b(b21to31), .out_c(matrixC21));
 processing_element_systolic_4x4_fp pe22(.reset(effective_rst), .clk(clk),  .in_a(a21to22), .in_b(b12to22), .out_a(a22to23), .out_b(b22to32), .out_c(matrixC22));
 processing_element_systolic_4x4_fp pe23(.reset(effective_rst), .clk(clk),  .in_a(a22to23), .in_b(b13to23), .out_a(a23to24), .out_b(b23to33), .out_c(matrixC23));

 processing_element_systolic_4x4_fp pe30(.reset(effective_rst), .clk(clk),  .in_a(a3),      .in_b(b20to30), .out_a(a30to31), .out_b(b30to40), .out_c(matrixC30));
 processing_element_systolic_4x4_fp pe31(.reset(effective_rst), .clk(clk),  .in_a(a30to31), .in_b(b21to31), .out_a(a31to32), .out_b(b31to41), .out_c(matrixC31));
 processing_element_systolic_4x4_fp pe32(.reset(effective_rst), .clk(clk),  .in_a(a31to32), .in_b(b22to32), .out_a(a32to33), .out_b(b32to42), .out_c(matrixC32));
 processing_element_systolic_4x4_fp pe33(.reset(effective_rst), .clk(clk),  .in_a(a32to33), .in_b(b23to33), .out_a(a33to34), .out_b(b33to43), .out_c(matrixC33));

assign a_data_out = {a33to34,a23to24,a13to14,a03to04};
assign b_data_out = {b33to43,b32to42,b31to41,b30to40};

endmodule



//////////////////////////////////////////////////////////////////////////
// Definition of a processing element (basically a MAC)
//////////////////////////////////////////////////////////////////////////
module  processing_element_systolic_4x4_fp(
 reset, 
 clk, 
 in_a,
 in_b, 
 out_a, 
 out_b, 
 out_c
 );

 input reset;
 input clk;
 input  [`DWIDTH-1:0] in_a;
 input  [`DWIDTH-1:0] in_b;
 output [`DWIDTH-1:0] out_a;
 output [`DWIDTH-1:0] out_b;
 output [`DWIDTH-1:0] out_c;  //reduced precision

 reg [`DWIDTH-1:0] out_a;
 reg [`DWIDTH-1:0] out_b;
 wire [`DWIDTH-1:0] out_c;

 wire [`DWIDTH-1:0] out_mac;

 assign out_c = out_mac;

 `ifdef complex_dsp
 mac_fp_16 u_mac(.a(in_a), .b(in_b), .out(out_mac), .reset(reset), .clk(clk));
 `else
 seq_mac_systolic_4x4_fp u_mac(.a(in_a), .b(in_b), .out(out_mac), .reset(reset), .clk(clk));
 `endif

 always @(posedge clk)begin
    if(reset) begin
      out_a<=0;
      out_b<=0;
    end
    else begin  
      out_a<=in_a;
      out_b<=in_b;
    end
 end
 
endmodule

//////////////////////////////////////////////////////////////////////////
// Multiply-and-accumulate (MAC) block
//////////////////////////////////////////////////////////////////////////
//module seq_mac_systolic_4x4_fp(a, b, out, reset, clk);
//input [`DWIDTH-1:0] a;
//input [`DWIDTH-1:0] b;
//input reset;
//input clk;
//output [`DWIDTH-1:0] out;
//
//reg [2*`DWIDTH-1:0] out_temp;
//wire [`DWIDTH-1:0] mul_out;
//wire [2*`DWIDTH-1:0] add_out;
//
//reg [`DWIDTH-1:0] a_flopped;
//reg [`DWIDTH-1:0] b_flopped;
//
//wire [2*`DWIDTH-1:0] mul_out_temp;
//reg [2*`DWIDTH-1:0] mul_out_temp_reg;
//
//always @(posedge clk) begin
//  if (reset) begin
//    a_flopped <= 0;
//    b_flopped <= 0;
//  end else begin
//    a_flopped <= a;
//    b_flopped <= b;
//  end
//end
//
////assign mul_out = a * b;
//qmult_systolic_4x4_fp mult_u1(.i_multiplicand(a_flopped), .i_multiplier(b_flopped), .o_result(mul_out_temp));
//
//always @(posedge clk) begin
//  if (reset) begin
//    mul_out_temp_reg <= 0;
//  end else begin
//    mul_out_temp_reg <= mul_out_temp;
//  end
//end
//
////we just truncate the higher bits of the product
////assign add_out = mul_out + out;
//qadd_systolic_4x4_fp add_u1(.a(out_temp), .b(mul_out_temp_reg), .c(add_out));
//
//always @(posedge clk) begin
//  if (reset) begin
//    out_temp <= 0;
//  end else begin
//    out_temp <= add_out;
//  end
//end
//
////down cast the result
//assign out = 
//    (out_temp[2*`DWIDTH-1] == 0) ?  //positive number
//        (
//           (|(out_temp[2*`DWIDTH-2 : `DWIDTH-1])) ?  //is any bit from 14:7 is 1, that means overlfow
//             {out_temp[2*`DWIDTH-1] , {(`DWIDTH-1){1'b1}}} : //sign bit and then all 1s
//             {out_temp[2*`DWIDTH-1] , out_temp[`DWIDTH-2:0]} 
//        )
//        : //negative number
//        (
//           (|(out_temp[2*`DWIDTH-2 : `DWIDTH-1])) ?  //is any bit from 14:7 is 0, that means overlfow
//             {out_temp[2*`DWIDTH-1] , out_temp[`DWIDTH-2:0]} :
//             {out_temp[2*`DWIDTH-1] , {(`DWIDTH-1){1'b0}}} //sign bit and then all 0s
//        );
//
//endmodule
//
//module qmult_systolic_4x4_fp(i_multiplicand,i_multiplier,o_result);
//input [`DWIDTH-1:0] i_multiplicand;
//input [`DWIDTH-1:0] i_multiplier;
//output [2*`DWIDTH-1:0] o_result;
//
//assign o_result = i_multiplicand * i_multiplier;
////DW02_mult #(`DWIDTH,`DWIDTH) u_mult(.A(i_multiplicand), .B(i_multiplier), .TC(1'b1), .PRODUCT(o_result));
//
//endmodule
//
//module qadd_systolic_4x4_fp(a,b,c);
//input [2*`DWIDTH-1:0] a;
//input [2*`DWIDTH-1:0] b;
//output [2*`DWIDTH-1:0] c;
//
//assign c = a + b;
////DW01_add #(`DWIDTH) u_add(.A(a), .B(b), .CI(1'b0), .SUM(c), .CO());
//endmodule

`ifndef complex_dsp

//////////////////////////////////////////////////////////////////////////
// Multiply-and-accumulate (MAC) block
//////////////////////////////////////////////////////////////////////////
module seq_mac_systolic_4x4_fp(a, b, out, reset, clk);
input [`DWIDTH-1:0] a;
input [`DWIDTH-1:0] b;
input reset;
input clk;
output [`DWIDTH-1:0] out;

reg [2*`DWIDTH-1:0] out_temp;
wire [2*`DWIDTH-1:0] mul_out;
wire [2*`DWIDTH-1:0] add_out;

reg [`DWIDTH-1:0] a_flopped;
reg [`DWIDTH-1:0] b_flopped;

wire [2*`DWIDTH-1:0] mul_out_temp;
reg [2*`DWIDTH-1:0] mul_out_temp_reg;

always @(posedge clk) begin
  if (reset) begin
    a_flopped <= 0;
    b_flopped <= 0;
  end else begin
    a_flopped <= a;
    b_flopped <= b;
  end
end

//assign mul_out = a * b;
qmult_systolic_4x4_fp mult_u1(.clk(clk), .rst(reset), .i_multiplicand(a_flopped), .i_multiplier(b_flopped), .o_result(mul_out_temp));

always @(posedge clk) begin
  if (reset) begin
    mul_out_temp_reg <= 0;
  end else begin
    mul_out_temp_reg <= mul_out_temp;
  end
end

assign mul_out = mul_out_temp_reg;

qadd_systolic_4x4_fp add_u1(.clk(clk), .rst(reset), .a(out_temp), .b(mul_out), .c(add_out));

always @(posedge clk) begin
  if (reset) begin
    out_temp <= 0;
  end else begin
    out_temp <= add_out;
  end
end

//fp32 to fp16 conversion
wire [15:0] fpadd_16_result;
fp32_to_fp16_systolic_4x4_fp u_32to16 (.a(out_temp), .b(out));

endmodule


//////////////////////////////////////////////////////////////////////////
// Multiplier
//////////////////////////////////////////////////////////////////////////
module qmult_systolic_4x4_fp(clk,rst,i_multiplicand,i_multiplier,o_result);
input clk;
input rst;
input [`DWIDTH-1:0] i_multiplicand;
input [`DWIDTH-1:0] i_multiplier;
output [2*`DWIDTH-1:0] o_result;

wire FPMult_16_systolic_4x4_fp_clk_NC;
wire FPMult_16_systolic_4x4_fp_rst_NC;
wire [15:0] FPMult_16_systolic_4x4_fp_result;
wire [4:0] FPMult_16_systolic_4x4_fp_flags;

FPMult_16_systolic_4x4_fp u_FPMult_16_systolic_4x4_fp(
   .clk(clk),
   .rst(rst),
   .a(i_multiplicand[15:0]),
   .b(i_multiplier[15:0]),
   .result(FPMult_16_systolic_4x4_fp_result),
   .flags(FPMult_16_systolic_4x4_fp_flags)
 );

//Convert fp16 to fp32
fp16_to_fp32_systolic_4x4_fp u_16to32 (.a(FPMult_16_systolic_4x4_fp_result), .b(o_result));

endmodule


//////////////////////////////////////////////////////////////////////////
// Adder
//////////////////////////////////////////////////////////////////////////
module qadd_systolic_4x4_fp(clk,rst,a,b,c);
input clk;
input rst;
input [2*`DWIDTH-1:0] a;
input [2*`DWIDTH-1:0] b;
output [2*`DWIDTH-1:0] c;

wire fpadd_32_clk_NC;
wire fpadd_32_rst_NC;
wire [4:0] fpadd_32_flags;

FPAddSub_single_systolic_4x4_fp u_fpaddsub_32(
  .clk(clk),
  .rst(rst),
  .a(a),
  .b(b),
  .operation(1'b0), 
  .result(c),
  .flags(fpadd_32_flags));

endmodule
`endif

`ifndef complex_dsp

//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////
// Definition of a 16-bit floating point multiplier
// This is a heavily modified version of:
// https://github.com/fbrosser/DSP48E1-FP/tree/master/src/FPMult
// Original author: Fredrik Brosser
// Abridged by: Samidh Mehta
//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////

module FPMult_16_systolic_4x4_fp(
		clk,
		rst,
		a,
		b,
		result,
		flags
    );
	
	// Input Ports
	input clk ;							// Clock
	input rst ;							// Reset signal
	input [`DWIDTH-1:0] a;						// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b;						// Input B, a 32-bit floating point number
	
	// Output ports
	output [`DWIDTH-1:0] result ;					// Product, result of the operation, 32-bit FP number
	output [4:0] flags ;						// Flags indicating exceptions according to IEEE754
	
	// Internal signals
	wire [`DWIDTH-1:0] Z_int ;					// Product, result of the operation, 32-bit FP number
	wire [4:0] Flags_int ;						// Flags indicating exceptions according to IEEE754
	
	wire Sa ;							// A's sign
	wire Sb ;							// B's sign
	wire Sp ;							// Product sign
	wire [`EXPONENT-1:0] Ea ;					// A's exponent
	wire [`EXPONENT-1:0] Eb ;					// B's exponent
	wire [2*`MANTISSA+1:0] Mp ;					// Product mantissa
	wire [4:0] InputExc ;						// Exceptions in inputs
	wire [`MANTISSA-1:0] NormM ;					// Normalized mantissa
	wire [`EXPONENT:0] NormE ;					// Normalized exponent
	wire [`MANTISSA:0] RoundM ;					// Normalized mantissa
	wire [`EXPONENT:0] RoundE ;					// Normalized exponent
	wire [`MANTISSA:0] RoundMP ;					// Normalized mantissa
	wire [`EXPONENT:0] RoundEP ;					// Normalized exponent
	wire GRS ;

	//reg [63:0] pipe_0;						// Pipeline register Input->Prep
	reg [2*`DWIDTH-1:0] pipe_0;					// Pipeline register Input->Prep

	//reg [92:0] pipe_1;						// Pipeline register Prep->Execute
	//reg [3*`MANTISSA+2*`EXPONENT+7:0] pipe_1;			// Pipeline register Prep->Execute
	reg [3*`MANTISSA+2*`EXPONENT+18:0] pipe_1;

	//reg [38:0] pipe_2;						// Pipeline register Execute->Normalize
	reg [`MANTISSA+`EXPONENT+7:0] pipe_2;				// Pipeline register Execute->Normalize
	
	//reg [72:0] pipe_3;						// Pipeline register Normalize->Round
	reg [2*`MANTISSA+2*`EXPONENT+10:0] pipe_3;			// Pipeline register Normalize->Round

	//reg [36:0] pipe_4;						// Pipeline register Round->Output
	reg [`DWIDTH+4:0] pipe_4;					// Pipeline register Round->Output
	
	assign result = pipe_4[`DWIDTH+4:5] ;
	assign flags = pipe_4[4:0] ;
	
	// Prepare the operands for alignment and check for exceptions
	FPMult_PrepModule_systolic_4x4_fp PrepModule(clk, rst, pipe_0[2*`DWIDTH-1:`DWIDTH], pipe_0[`DWIDTH-1:0], Sa, Sb, Ea[`EXPONENT-1:0], Eb[`EXPONENT-1:0], Mp[2*`MANTISSA+1:0], InputExc[4:0]) ;

	// Perform (unsigned) mantissa multiplication
	FPMult_ExecuteModule_systolic_4x4_fp ExecuteModule(pipe_1[3*`MANTISSA+`EXPONENT*2+7:2*`MANTISSA+2*`EXPONENT+8], pipe_1[2*`MANTISSA+2*`EXPONENT+7:2*`MANTISSA+7], pipe_1[2*`MANTISSA+6:5], pipe_1[2*`MANTISSA+2*`EXPONENT+6:2*`MANTISSA+`EXPONENT+7], pipe_1[2*`MANTISSA+`EXPONENT+6:2*`MANTISSA+7], pipe_1[2*`MANTISSA+2*`EXPONENT+8], pipe_1[2*`MANTISSA+2*`EXPONENT+7], Sp, NormE[`EXPONENT:0], NormM[`MANTISSA-1:0], GRS) ;

	// Round result and if necessary, perform a second (post-rounding) normalization step
	FPMult_NormalizeModule_systolic_4x4_fp NormalizeModule(pipe_2[`MANTISSA-1:0], pipe_2[`MANTISSA+`EXPONENT:`MANTISSA], RoundE[`EXPONENT:0], RoundEP[`EXPONENT:0], RoundM[`MANTISSA:0], RoundMP[`MANTISSA:0]) ;		

	// Round result and if necessary, perform a second (post-rounding) normalization step
	//FPMult_RoundModule_systolic_4x4_fp RoundModule(pipe_3[47:24], pipe_3[23:0], pipe_3[65:57], pipe_3[56:48], pipe_3[66], pipe_3[67], pipe_3[72:68], Z_int[31:0], Flags_int[4:0]) ;		
	FPMult_RoundModule_systolic_4x4_fp RoundModule(pipe_3[2*`MANTISSA+1:`MANTISSA+1], pipe_3[`MANTISSA:0], pipe_3[2*`MANTISSA+2*`EXPONENT+3:2*`MANTISSA+`EXPONENT+3], pipe_3[2*`MANTISSA+`EXPONENT+2:2*`MANTISSA+2], pipe_3[2*`MANTISSA+2*`EXPONENT+4], pipe_3[2*`MANTISSA+2*`EXPONENT+5], pipe_3[2*`MANTISSA+2*`EXPONENT+10:2*`MANTISSA+2*`EXPONENT+6], Z_int[`DWIDTH-1:0], Flags_int[4:0]) ;		

//adding always@ (*) instead of posedge clock to make design combinational
	always @ (posedge clk) begin	
		if(rst) begin
			pipe_0 <= 0;
			pipe_1 <= 0;
			pipe_2 <= 0; 
			pipe_3 <= 0;
			pipe_4 <= 0;
		end 
		else begin		
			/* PIPE 0
				[2*`DWIDTH-1:`DWIDTH] A
				[`DWIDTH-1:0] B
			*/
                       pipe_0 <= {a, b} ;


			/* PIPE 1
				[2*`EXPONENT+3*`MANTISSA + 18: 2*`EXPONENT+2*`MANTISSA + 18] //pipe_0[`DWIDTH+`MANTISSA-1:`DWIDTH] , mantissa of A
				[2*`EXPONENT+2*`MANTISSA + 17 :2*`EXPONENT+2*`MANTISSA + 9] // pipe_0[8:0]
				[2*`EXPONENT+2*`MANTISSA + 8] Sa
				[2*`EXPONENT+2*`MANTISSA + 7] Sb
				[2*`EXPONENT+2*`MANTISSA + 6:`EXPONENT+2*`MANTISSA+7] Ea
				[`EXPONENT +2*`MANTISSA+6:2*`MANTISSA+7] Eb
				[2*`MANTISSA+1+5:5] Mp
				[4:0] InputExc
			*/
			//pipe_1 <= {pipe_0[`DWIDTH+`MANTISSA-1:`DWIDTH], pipe_0[`MANTISSA_MUL_SPLIT_LSB-1:0], Sa, Sb, Ea[`EXPONENT-1:0], Eb[`EXPONENT-1:0], Mp[2*`MANTISSA-1:0], InputExc[4:0]} ;
			pipe_1 <= {pipe_0[`DWIDTH+`MANTISSA-1:`DWIDTH], pipe_0[8:0], Sa, Sb, Ea[`EXPONENT-1:0], Eb[`EXPONENT-1:0], Mp[2*`MANTISSA+1:0], InputExc[4:0]} ;
			
			/* PIPE 2
				[`EXPONENT + `MANTISSA + 7:`EXPONENT + `MANTISSA + 3] InputExc
				[`EXPONENT + `MANTISSA + 2] GRS
				[`EXPONENT + `MANTISSA + 1] Sp
				[`EXPONENT + `MANTISSA:`MANTISSA] NormE
				[`MANTISSA-1:0] NormM
			*/
			pipe_2 <= {pipe_1[4:0], GRS, Sp, NormE[`EXPONENT:0], NormM[`MANTISSA-1:0]} ;
			/* PIPE 3
				[2*`EXPONENT+2*`MANTISSA+10:2*`EXPONENT+2*`MANTISSA+6] InputExc
				[2*`EXPONENT+2*`MANTISSA+5] GRS
				[2*`EXPONENT+2*`MANTISSA+4] Sp	
				[2*`EXPONENT+2*`MANTISSA+3:`EXPONENT+2*`MANTISSA+3] RoundE
				[`EXPONENT+2*`MANTISSA+2:2*`MANTISSA+2] RoundEP
				[2*`MANTISSA+1:`MANTISSA+1] RoundM
				[`MANTISSA:0] RoundMP
			*/
			pipe_3 <= {pipe_2[`EXPONENT+`MANTISSA+7:`EXPONENT+`MANTISSA+1], RoundE[`EXPONENT:0], RoundEP[`EXPONENT:0], RoundM[`MANTISSA:0], RoundMP[`MANTISSA:0]} ;
			/* PIPE 4
				[`DWIDTH+4:5] Z
				[4:0] Flags
			*/				
			pipe_4 <= {Z_int[`DWIDTH-1:0], Flags_int[4:0]} ;
		end
	end
		
endmodule



module FPMult_PrepModule_systolic_4x4_fp (
		clk,
		rst,
		a,
		b,
		Sa,
		Sb,
		Ea,
		Eb,
		Mp,
		InputExc
	);
	
	// Input ports
	input clk ;
	input rst ;
	input [`DWIDTH-1:0] a ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b ;								// Input B, a 32-bit floating point number
	
	// Output ports
	output Sa ;										// A's sign
	output Sb ;										// B's sign
	output [`EXPONENT-1:0] Ea ;								// A's exponent
	output [`EXPONENT-1:0] Eb ;								// B's exponent
	output [2*`MANTISSA+1:0] Mp ;							// Mantissa product
	output [4:0] InputExc ;						// Input numbers are exceptions
	
	// Internal signals							// If signal is high...
	wire ANaN ;										// A is a signalling NaN
	wire BNaN ;										// B is a signalling NaN
	wire AInf ;										// A is infinity
	wire BInf ;										// B is infinity
    wire [`MANTISSA-1:0] Ma;
    wire [`MANTISSA-1:0] Mb;
	
	assign ANaN = &(a[`DWIDTH-2:`MANTISSA]) &  |(a[`DWIDTH-2:`MANTISSA]) ;			// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(b[`DWIDTH-2:`MANTISSA]) &  |(b[`MANTISSA-1:0]);			// All one exponent and not all zero mantissa - NaN
	assign AInf = &(a[`DWIDTH-2:`MANTISSA]) & ~|(a[`DWIDTH-2:`MANTISSA]) ;		// All one exponent and all zero mantissa - Infinity
	assign BInf = &(b[`DWIDTH-2:`MANTISSA]) & ~|(b[`DWIDTH-2:`MANTISSA]) ;		// All one exponent and all zero mantissa - Infinity
	
	// Check for any exceptions and put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	//assign InputExc = {(ANaN | ANaN | BNaN |BNaN), ANaN, ANaN, BNaN,BNaN} ;
	
	// Take input numbers apart
	assign Sa = a[`DWIDTH-1] ;							// A's sign
	assign Sb = b[`DWIDTH-1] ;							// B's sign
	assign Ea = a[`DWIDTH-2:`MANTISSA];						// Store A's exponent in Ea, unless A is an exception
	assign Eb = b[`DWIDTH-2:`MANTISSA];						// Store B's exponent in Eb, unless B is an exception	
//    assign Ma = a[`MANTISSA_MSB:`MANTISSA_LSB];
  //  assign Mb = b[`MANTISSA_MSB:`MANTISSA_LSB];
	


	//assign Mp = ({4'b0001, a[`MANTISSA-1:0]}*{4'b0001, b[`MANTISSA-1:9]}) ;
	assign Mp = ({1'b1,a[`MANTISSA-1:0]}*{1'b1, b[`MANTISSA-1:0]}) ;

	
    //We multiply part of the mantissa here
    //Full mantissa of A
    //Bits MANTISSA_MUL_SPLIT_MSB:MANTISSA_MUL_SPLIT_LSB of B
   // wire [`ACTUAL_MANTISSA-1:0] inp_A;
   // wire [`ACTUAL_MANTISSA-1:0] inp_B;
   // assign inp_A = {1'b1, Ma};
   // assign inp_B = {{(`MANTISSA-(`MANTISSA_MUL_SPLIT_MSB-`MANTISSA_MUL_SPLIT_LSB+1)){1'b0}}, 1'b1, Mb[`MANTISSA_MUL_SPLIT_MSB:`MANTISSA_MUL_SPLIT_LSB]};
   // DW02_mult #(`ACTUAL_MANTISSA,`ACTUAL_MANTISSA) u_mult(.A(inp_A), .B(inp_B), .TC(1'b0), .PRODUCT(Mp));
endmodule


module FPMult_ExecuteModule_systolic_4x4_fp(
		a,
		b,
		MpC,
		Ea,
		Eb,
		Sa,
		Sb,
		Sp,
		NormE,
		NormM,
		GRS
    );

	// Input ports
	input [`MANTISSA-1:0] a ;
	input [2*`EXPONENT:0] b ;
	input [2*`MANTISSA+1:0] MpC ;
	input [`EXPONENT-1:0] Ea ;						// A's exponent
	input [`EXPONENT-1:0] Eb ;						// B's exponent
	input Sa ;								// A's sign
	input Sb ;								// B's sign
	
	// Output ports
	output Sp ;								// Product sign
	output [`EXPONENT:0] NormE ;													// Normalized exponent
	output [`MANTISSA-1:0] NormM ;												// Normalized mantissa
	output GRS ;
	
	wire [2*`MANTISSA+1:0] Mp ;
	
	assign Sp = (Sa ^ Sb) ;												// Equal signs give a positive product
	
   // wire [`ACTUAL_MANTISSA-1:0] inp_a;
   // wire [`ACTUAL_MANTISSA-1:0] inp_b;
   // assign inp_a = {1'b1, a};
   // assign inp_b = {{(`MANTISSA-`MANTISSA_MUL_SPLIT_LSB){1'b0}}, 1'b0, b};
   // DW02_mult #(`ACTUAL_MANTISSA,`ACTUAL_MANTISSA) u_mult(.A(inp_a), .B(inp_b), .TC(1'b0), .PRODUCT(Mp_temp));
   // DW01_add #(2*`ACTUAL_MANTISSA) u_add(.A(Mp_temp), .B(MpC<<`MANTISSA_MUL_SPLIT_LSB), .CI(1'b0), .SUM(Mp), .CO());

	//assign Mp = (MpC<<(2*`EXPONENT+1)) + ({4'b0001, a[`MANTISSA-1:0]}*{1'b0, b[2*`EXPONENT:0]}) ;
	assign Mp = MpC;


	assign NormM = (Mp[2*`MANTISSA+1] ? Mp[2*`MANTISSA:`MANTISSA+1] : Mp[2*`MANTISSA-1:`MANTISSA]); 	// Check for overflow
	assign NormE = (Ea + Eb + Mp[2*`MANTISSA+1]);								// If so, increment exponent
	
	assign GRS = ((Mp[`MANTISSA]&(Mp[`MANTISSA+1]))|(|Mp[`MANTISSA-1:0])) ;
	
endmodule

module FPMult_NormalizeModule_systolic_4x4_fp(
		NormM,
		NormE,
		RoundE,
		RoundEP,
		RoundM,
		RoundMP
    );

	// Input Ports
	input [`MANTISSA-1:0] NormM ;									// Normalized mantissa
	input [`EXPONENT:0] NormE ;									// Normalized exponent

	// Output Ports
	output [`EXPONENT:0] RoundE ;
	output [`EXPONENT:0] RoundEP ;
	output [`MANTISSA:0] RoundM ;
	output [`MANTISSA:0] RoundMP ; 
	
// EXPONENT = 5 
// EXPONENT -1 = 4
// NEED to subtract 2^4 -1 = 15

wire [`EXPONENT-1 : 0] bias;

assign bias =  ((1<< (`EXPONENT -1)) -1);

	assign RoundE = NormE - bias ;
	assign RoundEP = NormE - bias -1 ;
	assign RoundM = NormM ;
	assign RoundMP = NormM ;

endmodule

module FPMult_RoundModule_systolic_4x4_fp(
		RoundM,
		RoundMP,
		RoundE,
		RoundEP,
		Sp,
		GRS,
		InputExc,
		Z,
		Flags
    );

	// Input Ports
	input [`MANTISSA:0] RoundM ;									// Normalized mantissa
	input [`MANTISSA:0] RoundMP ;									// Normalized exponent
	input [`EXPONENT:0] RoundE ;									// Normalized mantissa + 1
	input [`EXPONENT:0] RoundEP ;									// Normalized exponent + 1
	input Sp ;												// Product sign
	input GRS ;
	input [4:0] InputExc ;
	
	// Output Ports
	output [`DWIDTH-1:0] Z ;										// Final product
	output [4:0] Flags ;
	
	// Internal Signals
	wire [`EXPONENT:0] FinalE ;									// Rounded exponent
	wire [`MANTISSA:0] FinalM;
	wire [`MANTISSA:0] PreShiftM;
	
	assign PreShiftM = GRS ? RoundMP : RoundM ;	// Round up if R and (G or S)
	
	// Post rounding normalization (potential one bit shift> use shifted mantissa if there is overflow)
	assign FinalM = (PreShiftM[`MANTISSA] ? {1'b0, PreShiftM[`MANTISSA:1]} : PreShiftM[`MANTISSA:0]) ;
	
	assign FinalE = (PreShiftM[`MANTISSA] ? RoundEP : RoundE) ; // Increment exponent if a shift was done
	
	assign Z = {Sp, FinalE[`EXPONENT-1:0], FinalM[`MANTISSA-1:0]} ;   // Putting the pieces together
	assign Flags = InputExc[4:0];

endmodule

`endif

 
//////////////////////////////////////////////////////////////////////////
// A floating point 16-bit to floating point 32-bit converter
//////////////////////////////////////////////////////////////////////////
`ifndef complex_dsp
module fp16_to_fp32_systolic_4x4_fp (input [15:0] a , output [31:0] b);

reg [31:0]b_temp;
reg [3:0] j;
reg [3:0] k;
reg [3:0] k_temp;
always @ (*) begin

if ( a [14: 0] == 15'b0 ) begin //signed zero
	b_temp [31] = a[15]; //sign bit
	b_temp[30:0] = 31'b0;
end

else begin

	if ( a[14 : 10] == 5'b0 ) begin //denormalized (covert to normalized)
		
		for (j=0; j<=9; j=j+1) begin
			if (a[j] == 1'b1) begin 
			    k_temp = j;	
			end
		end
	k = 9 - k_temp;

	b_temp [22:0] = ( (a [9:0] << (k+1'b1)) & 10'h3FF ) << 13;
	b_temp [30:23] =  7'd127 - 4'd15 - k;
	b_temp [31] = a[15];
	end

	else if ( a[14 : 10] == 5'b11111 ) begin //Infinity/ NAN
	b_temp [22:0] = a [9:0] << 13;
	b_temp [30:23] = 8'hFF;
	b_temp [31] = a[15];
	end

	else begin //Normalized Number
	b_temp [22:0] = a [9:0] << 13;
	b_temp [30:23] =  7'd127 - 4'd15 + a[14:10];
	b_temp [31] = a[15];
	end
end
end

assign b = b_temp;


endmodule

//////////////////////////////////////////////////////////////////////////
// A floating point 32-bit to floating point 16-bit converter
//////////////////////////////////////////////////////////////////////////
module fp32_to_fp16_systolic_4x4_fp (input [31:0] a , output [15:0] b);

reg [15:0]b_temp;
//integer j;
//reg [3:0]k;
always @ (*) begin

if ( a [30: 0] == 15'b0 ) begin //signed zero
	b_temp [15] = a[30]; //sign bit
	b_temp [14:0] = 15'b0; 
end

else begin

	if ( a[30 : 23] <= 8'd112  &&  a[30 : 23] >= 8'd103 ) begin //denormalized (covert to normalized)
		
	b_temp [9:0] = {1'b1, a[22:13]} >> {8'd112 - a[30 : 23] + 1'b1} ;  
	b_temp [14:10] =  5'b0;
	b_temp [15] = a[31];
	end

	else if ( a[ 30 : 23] == 8'b11111111 ) begin //Infinity/ NAN
	b_temp [9:0] = a [22:13];
	b_temp [14:10] = 5'h1F;
	b_temp [15] = a[31];
	end

	else begin //Normalized Number
	b_temp [9:0] = a [22:13];
	b_temp [14:10] = 4'd15 - 7'd127  + a[30:23]; //number should be in the range which can be depicted by fp16 (exp for fp32: 70h, 8Eh ; normalized exp for fp32: -15 to 15)
	b_temp [15] = a[31];
	end
end
end

assign b = b_temp;


endmodule
`endif

//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////
// Definition of a 32-bit floating point adder/subtractor
// This is a heavily modified version of:
// https://github.com/fbrosser/DSP48E1-FP/tree/master/src/FP_AddSub
// Original author: Fredrik Brosser
// Abridged by: Samidh Mehta
//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////

`ifndef complex_dsp
module FPAddSub_single_systolic_4x4_fp(
		clk,
		rst,
		a,
		b,
		operation,
		result,
		flags
	);

// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [31:0] a ;								// Input A, a 32-bit floating point number
	input [31:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [31:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754

	reg [68:0]pipe_1;
	reg [54:0]pipe_2;
	reg [45:0]pipe_3;


//internal module wires

//output ports
	wire Opout;
	wire Sa;
	wire Sb;
	wire MaxAB;
	wire [7:0] CExp;
	wire [4:0] Shift;
	wire [22:0] Mmax;
	wire [4:0] InputExc;
	wire [23:0] Mmin_3;

	wire [32:0] SumS_5 ;
	wire [4:0] Shift_1;							
	wire PSgn ;							
	wire Opr ;	
	
	wire [22:0] NormM ;				// Normalized mantissa
	wire [8:0] NormE ;					// Adjusted exponent
	wire ZeroSum ;						// Zero flag
	wire NegE ;							// Flag indicating negative exponent
	wire R ;								// Round bit
	wire S ;								// Final sticky bit
	wire FG ;

FPAddSub_a_systolic_4x4_fp M1(a,b,operation,Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3);

FPAddSub_b_systolic_4x4_fp M2(pipe_1[51:29],pipe_1[23:0],pipe_1[67],pipe_1[66],pipe_1[65],pipe_1[68],SumS_5,Shift_1,PSgn,Opr);

FPAddSub_c_systolic_4x4_fp M3(pipe_2[54:22],pipe_2[21:17],pipe_2[16:9],NormM,NormE,ZeroSum,NegE,R,S,FG);

FPAddSub_d_systolic_4x4_fp M4(pipe_3[13],pipe_3[22:14],pipe_3[45:23],pipe_3[11],pipe_3[10],pipe_3[9],pipe_3[8],pipe_3[7],pipe_3[6],pipe_3[5],pipe_3[12],pipe_3[4:0],result,flags );


always @ (posedge clk) begin	
		if(rst) begin
			pipe_1 <= 0;
			pipe_2 <= 0;
			pipe_3 <= 0;
		end 
		else begin
/*
pipe_1:
	[68] Opout;
	[67] Sa;
	[66] Sb;
	[65] MaxAB;
	[64:57] CExp;
	[56:52] Shift;
	[51:29] Mmax;
	[28:24] InputExc;
	[23:0] Mmin_3;	
*/

pipe_1 <= {Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3};

/*
pipe_2:
	[54:22]SumS_5;
	[21:17]Shift;
	[16:9]CExp;	
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_2 <= {SumS_5,Shift_1,pipe_1[64:57], pipe_1[67], pipe_1[66], pipe_1[68], pipe_1[65], pipe_1[28:24] };

/*
pipe_3:
	[45:23] NormM ;				
	[22:14] NormE ;					
	[13]ZeroSum ;						
	[12]NegE ;							
	[11]R ;								
	[10]S ;								
	[9]FG ;
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_3 <= {NormM,NormE,ZeroSum,NegE,R,S,FG, pipe_2[8], pipe_2[7], pipe_2[6], pipe_2[5], pipe_2[4:0] };

end
end

endmodule

// Prealign + Align + Shift 1 + Shift 2
module FPAddSub_a_systolic_4x4_fp(
		A,
		B,
		operation,
		Opout,
		Sa,
		Sb,
		MaxAB,
		CExp,
		Shift,
		Mmax,
		InputExc,
		Mmin_3
		
		
	);
	
	// Input ports
	input [31:0] A ;										// Input A, a 32-bit floating point number
	input [31:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	//output ports
	output Opout;
	output Sa;
	output Sb;
	output MaxAB;
	output [7:0] CExp;
	output [4:0] Shift;
	output [22:0] Mmax;
	output [4:0] InputExc;
	output [23:0] Mmin_3;	
							
	wire [9:0] ShiftDet ;							
	wire [30:0] Aout ;
	wire [30:0] Bout ;
	

	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [7:0] DAB ;										// ExpA - ExpB					
	wire [7:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[30:23]) & |(A[22:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[30:23]) & |(B[22:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[30:23]) & ~|(A[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[30:23]) & ~|(B[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
  assign DAB = (A[30:23] + ~(B[30:23]) + 1) ;
	assign DBA = (B[30:23] + ~(A[30:23]) + 1) ;

	assign Sa = A[31] ;									// A's sign bit
	assign Sb = B[31] ;									// B's sign	bit
	assign ShiftDet = {DBA[4:0], DAB[4:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[30:0] ;
	assign Bout = B[30:0] ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Output ports
													// Number of steps to smaller mantissa shift right
	wire [22:0] Mmin_1 ;							// Smaller mantissa 
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (Aout[30:0] < Bout[30:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[9:5] : ShiftDet[4:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin_1 = MaxAB ? Aout[22:0] : Bout[22:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? Bout[22:0]: Aout[22:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? Bout[30:23] : Aout[30:23]) ;	

// Input ports
					// Smaller mantissa after 16|12|8|4 shift
	wire [2:0] Shift_1 ;						// Shift amount
	
	assign Shift_1 = Shift [4:2];

	wire [23:0] Mmin_2 ;						// The smaller mantissa
	
	// Internal signals
	reg	  [23:0]		Lvl1;
	reg	  [23:0]		Lvl2;
	wire    [47:0]    Stage1;	
	integer           i;                // Loop variable
	
	always @(*) begin						
		// Rotate by 16?
		Lvl1 <= Shift_1[2] ? {17'b00000000000000001, Mmin_1[22:16]} : {1'b1, Mmin_1}; 
	end
	
	assign Stage1 = {Lvl1, Lvl1};
	
	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift_1[1:0])
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[23:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[23:19] <= 0; end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end Lvl2[23:15] <= 0; end
			// Rotate by 12	
			2'b11:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[23:11] <= 0; end
	  endcase
	end
	
	// Assign output to next shift stage
	assign Mmin_2 = Lvl2;
								// Smaller mantissa after 16|12|8|4 shift
	wire [1:0] Shift_2 ;						// Shift amount
	
	assign Shift_2 =Shift  [1:0] ;
					// The smaller mantissa
	
	// Internal Signal
	reg	  [23:0]		Lvl3;
	wire    [47:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {Mmin_2, Mmin_2};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_2[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[23:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end Lvl3[23] <= 0; end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end Lvl3[23:22] <= 0; end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end Lvl3[23:21] <= 0; end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin_3 = Lvl3;	

	
endmodule

module FPAddSub_b_systolic_4x4_fp(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		SumS_5,
		Shift,
		PSgn,
		Opr
);
	input [22:0] Mmax ;					// The larger mantissa
	input [23:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	wire [32:0] Sum ;	
						// Output ports
	output [32:0] SumS_5 ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount				// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation

	// Perform effective operation
	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, 8'b00000000} - {Mmin, 8'b00000000}) : ({1'b1, Mmax, 8'b00000000} + {Mmin, 8'b00000000}) ;
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

		// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[32] ? 5'b00000 :	 
		Sum[31] ? 5'b00001 : 
		Sum[30] ? 5'b00010 : 
		Sum[29] ? 5'b00011 : 
		Sum[28] ? 5'b00100 : 
		Sum[27] ? 5'b00101 : 
		Sum[26] ? 5'b00110 : 
		Sum[25] ? 5'b00111 :
		Sum[24] ? 5'b01000 :
		Sum[23] ? 5'b01001 :
		Sum[22] ? 5'b01010 :
		Sum[21] ? 5'b01011 :
		Sum[20] ? 5'b01100 :
		Sum[19] ? 5'b01101 :
		Sum[18] ? 5'b01110 :
		Sum[17] ? 5'b01111 :
		Sum[16] ? 5'b10000 :
		Sum[15] ? 5'b10001 :
		Sum[14] ? 5'b10010 :
		Sum[13] ? 5'b10011 :
		Sum[12] ? 5'b10100 :
		Sum[11] ? 5'b10101 :
		Sum[10] ? 5'b10110 :
		Sum[9] ? 5'b10111 :
		Sum[8] ? 5'b11000 :
		Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [32:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[16:0], 16'b0000000000000000} : Sum; 
	end
	
	// Assign outputs
	assign SumS_5 = Lvl1;	

endmodule

module FPAddSub_c_systolic_4x4_fp(
		SumS_5,
		Shift,
		CExp,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [32:0] SumS_5 ;						// Smaller mantissa after 16|12|8|4 shift
	
	input [4:0] Shift ;						// Shift amount
	
// Input ports
	
	input [7:0] CExp ;
	

	// Output ports
	output [22:0] NormM ;				// Normalized mantissa
	output [8:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;


	wire [3:0]Shift_1;
	assign Shift_1 = Shift [3:0];
	// Output ports
	wire [32:0] SumS_7 ;						// The smaller mantissa
	
	reg	  [32:0]		Lvl2;
	wire    [65:0]    Stage1;	
	reg	  [32:0]		Lvl3;
	wire    [65:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {SumS_5, SumS_5};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: Lvl2 <= Stage1[32:0];       		
			// Rotate by 4
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
			// Rotate by 8
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
			// Rotate by 12
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_1[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[32:0];
			// Rotate by 1
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
			// Rotate by 2
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
			// Rotate by 3
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
	  endcase
	end
	
	// Assign outputs
	assign SumS_7 = Lvl3;						// Take out smaller mantissa



	
	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [8:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [8:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = SumS_7[32] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|SumS_7 ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[8] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = SumS_7[31:9] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = SumS_7[8] ; 
	assign R = SumS_7[7] ;
	assign S = |SumS_7[6:0] ;		
	
endmodule

module FPAddSub_d_systolic_4x4_fp(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		NegE,
		InputExc,
		P,
		Flags 
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [8:0] NormE ;				// Normalized exponent
	input [22:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	

	input NegE ;						// Negative exponent?
	input [4:0] InputExc ;					// Exceptions in inputs A and B

	// Output ports
	output [31:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// 
	wire [31:0] Z ;					// Final result
	wire EOF ;
	
	// Internal signals
	wire [23:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [22:0] RoundM ;				// The final rounded sum
	wire [8:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	wire FSgn;
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[22:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[23] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? 8'b00000000 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[7:0], RoundM[22:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[8];

/////////////////////////////////////////////////////////////////////////////////////////////////////////



	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[30:23]) & ~|(Z[30:23]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule
`endif

module dbram_2048_60bit (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b,reset
); 

parameter AWIDTH=11;
parameter NUM_WORDS=2048;
parameter DWIDTH=60;
input clk, reset;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

reg count; 

always@(posedge clk) begin 

if (reset) begin 
	count <= 1'b0; 
end
else begin 
	count <= ~count; 
end

end

wire [(AWIDTH-1):0] address_a1,address_a2;
wire [(AWIDTH-1):0] address_b1,address_b2;
wire  wren_a1,wren_a2;
wire  wren_b1,wren_b2;
wire [(DWIDTH-1):0] data_a1,data_a2;
wire [(DWIDTH-1):0] data_b1,data_b2;
wire [(DWIDTH-1):0] out_a1,out_a2;
wire [(DWIDTH-1):0] out_b1,out_b2;

assign address_a1 = count|address_a; 
assign address_a2 = (~count)|address_a;
assign address_b1 = count|address_b; 
assign address_b2 = (~count)|address_b;
assign wren_a1 = count|wren_a; 
assign wren_a2 = (~count)|wren_a; 
assign wren_b1 = count|wren_b; 
assign wren_b2 = (~count)|wren_b; 
assign data_a1 = count|data_a;
assign data_a2 = (~count)|data_a;
assign data_b1 = count|data_b;
assign data_b2 = (~count)|data_b;
always@(posedge clk) begin
out_a <= count?out_a1:out_a2;
out_b <= count?out_b1:out_b2;
end

dpram_2048_60bit_db inst1(.clk(clk),.address_a(address_a1),.address_b(address_b1),.wren_a(wren_a1),.wren_b(wren_b1),.data_a(data_a1),.data_b(data_b1),.out_a(out_a1),.out_b(out_b1));
dpram_2048_60bit_db inst2(.clk(clk),.address_a(address_a2),.address_b(address_b2),.wren_a(wren_a2),.wren_b(wren_b2),.data_a(data_a2),.data_b(data_b2),.out_a(out_a2),.out_b(out_b2));


endmodule

module dpram_2048_60bit_db (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b
);
parameter AWIDTH=11;
parameter NUM_WORDS=2048;
parameter DWIDTH=60;
input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren_a) 
      ram[address_a] <= data_a;
  if (wren_b) 
      ram[address_b] <= data_b;

  out_a <= ram[address_a];
  out_b <= ram[address_b];
end
  

`else

defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

dual_port_ram u_dual_port_ram(
.addr1(address_a),
.we1(wren_a),
.data1(data_a),
.out1(out_a),
.addr2(address_b),
.we2(wren_b),
.data2(data_b),
.out2(out_b),
.clk(clk)
);

`endif
endmodule
module dbram_4096_40bit (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b,reset
); 

parameter AWIDTH=12;
parameter NUM_WORDS=4096;
parameter DWIDTH=40;
input clk, reset;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

reg count; 

always@(posedge clk) begin 

if (reset) begin 
	count <= 1'b0; 
end
else begin 
	count <= ~count; 
end

end

wire [(AWIDTH-1):0] address_a1,address_a2;
wire [(AWIDTH-1):0] address_b1,address_b2;
wire  wren_a1,wren_a2;
wire  wren_b1,wren_b2;
wire [(DWIDTH-1):0] data_a1,data_a2;
wire [(DWIDTH-1):0] data_b1,data_b2;
wire [(DWIDTH-1):0] out_a1,out_a2;
wire [(DWIDTH-1):0] out_b1,out_b2;

assign address_a1 = count|address_a; 
assign address_a2 = (~count)|address_a;
assign address_b1 = count|address_b; 
assign address_b2 = (~count)|address_b;
assign wren_a1 = count|wren_a; 
assign wren_a2 = (~count)|wren_a; 
assign wren_b1 = count|wren_b; 
assign wren_b2 = (~count)|wren_b; 
assign data_a1 = count|data_a;
assign data_a2 = (~count)|data_a;
assign data_b1 = count|data_b;
assign data_b2 = (~count)|data_b;
always@(posedge clk) begin
out_a <= count?out_a1:out_a2;
out_b <= count?out_b1:out_b2;
end
dpram_4096_40bit_db inst1(.clk(clk),.address_a(address_a1),.address_b(address_b1),.wren_a(wren_a1),.wren_b(wren_b1),.data_a(data_a1),.data_b(data_b1),.out_a(out_a1),.out_b(out_b1));
dpram_4096_40bit_db inst2(.clk(clk),.address_a(address_a2),.address_b(address_b2),.wren_a(wren_a2),.wren_b(wren_b2),.data_a(data_a2),.data_b(data_b2),.out_a(out_a2),.out_b(out_b2));


endmodule

module dpram_4096_40bit_db (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b
);
parameter AWIDTH=12;
parameter NUM_WORDS=4096;
parameter DWIDTH=40;
input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren_a) 
      ram[address_a] <= data_a;
  if (wren_b) 
      ram[address_b] <= data_b;
  
  out_a <= ram[address_a];
  out_b <= ram[address_b];
end

`else

defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

dual_port_ram u_dual_port_ram(
.addr1(address_a),
.we1(wren_a),
.data1(data_a),
.out1(out_a),
.addr2(address_b),
.we2(wren_b),
.data2(data_b),
.out2(out_b),
.clk(clk)
);

`endif
endmodule
module dbram_4096_60bit (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b,reset
); 

parameter AWIDTH=12;
parameter NUM_WORDS=4096;
parameter DWIDTH=60;
input clk,reset;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

reg count; 

always@(posedge clk) begin 

if (reset) begin 
	count <= 1'b0; 
end
else begin 
	count <= ~count; 
end

end

wire [(AWIDTH-1):0] address_a1,address_a2;
wire [(AWIDTH-1):0] address_b1,address_b2;
wire  wren_a1,wren_a2;
wire  wren_b1,wren_b2;
wire [(DWIDTH-1):0] data_a1,data_a2;
wire [(DWIDTH-1):0] data_b1,data_b2;
wire [(DWIDTH-1):0] out_a1,out_a2;
wire [(DWIDTH-1):0] out_b1,out_b2;

assign address_a1 = count|address_a; 
assign address_a2 = (~count)|address_a;
assign address_b1 = count|address_b; 
assign address_b2 = (~count)|address_b;
assign wren_a1 = count|wren_a; 
assign wren_a2 = (~count)|wren_a; 
assign wren_b1 = count|wren_b; 
assign wren_b2 = (~count)|wren_b; 
assign data_a1 = count|data_a;
assign data_a2 = (~count)|data_a;
assign data_b1 = count|data_b;
assign data_b2 = (~count)|data_b;
always@(posedge clk) begin
out_a <= count?out_a1:out_a2;
out_b <= count?out_b1:out_b2;
end

dpram_4096_60bit_db inst1(.clk(clk),.address_a(address_a1),.address_b(address_b1),.wren_a(wren_a1),.wren_b(wren_b1),.data_a(data_a1),.data_b(data_b1),.out_a(out_a1),.out_b(out_b1));
dpram_4096_60bit_db inst2(.clk(clk),.address_a(address_a2),.address_b(address_b2),.wren_a(wren_a2),.wren_b(wren_b2),.data_a(data_a2),.data_b(data_b2),.out_a(out_a2),.out_b(out_b2));


endmodule

module dpram_4096_60bit_db (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b
);
parameter AWIDTH=12;
parameter NUM_WORDS=4096;
parameter DWIDTH=60;
input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren_a) 
      ram[address_a] <= data_a;
  if (wren_b) 
      ram[address_b] <= data_b;
      
  out_a <= ram[address_a];
  out_b <= ram[address_b];
end

`else
defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

dual_port_ram u_dual_port_ram(
.addr1(address_a),
.we1(wren_a),
.data1(data_a),
.out1(out_a),
.addr2(address_b),
.we2(wren_b),
.data2(data_b),
.out2(out_b),
.clk(clk)
);

`endif
endmodule
`define DWIDTH 16
`define DESIGN_SIZE 32
`define MASK_WIDTH 2

module activation_32_16bit(
    input activation_type,
    input enable_activation,
    input in_data_available,
    input [`DESIGN_SIZE*`DWIDTH-1:0] inp_data,
    output [`DESIGN_SIZE*`DWIDTH-1:0] out_data,
    output out_data_available,
    input [`MASK_WIDTH-1:0] validity_mask,
    output done_activation,
    input clk,
    input reset
);

reg  done_activation_internal;
reg  out_data_available_internal;
wire [`DESIGN_SIZE*`DWIDTH-1:0] out_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] slope_applied_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] intercept_applied_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] relu_applied_data_internal;
reg [31:0] i;
reg [31:0] cycle_count;
reg activation_in_progress;

reg [(`DESIGN_SIZE*4)-1:0] address;
reg [(`DESIGN_SIZE*8)-1:0] data_slope;
reg [(`DESIGN_SIZE*8)-1:0] data_slope_flopped;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept_delayed;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept_flopped;

reg in_data_available_flopped;
reg [`DESIGN_SIZE*`DWIDTH-1:0] inp_data_flopped;

always @(posedge clk) begin
  if (reset) begin
    inp_data_flopped <= 0;
    data_slope_flopped <= 0;
  end else begin
    inp_data_flopped <= inp_data;
    data_slope_flopped <= data_slope;
  end
end

// If the activation block is not enabled, just forward the input data
assign out_data             = enable_activation ? out_data_internal : inp_data_flopped;
assign done_activation      = enable_activation ? done_activation_internal : 1'b1;
assign out_data_available   = enable_activation ? out_data_available_internal : in_data_available_flopped;

always @(posedge clk) begin
   if (reset || ~enable_activation) begin
      slope_applied_data_internal     <= 0;
      intercept_applied_data_internal <= 0; 
      relu_applied_data_internal      <= 0; 
      data_intercept_delayed      <= 0;
      data_intercept_flopped      <= 0;
      done_activation_internal    <= 0;
      out_data_available_internal <= 0;
      cycle_count                 <= 0;
      activation_in_progress      <= 0;
      in_data_available_flopped <= in_data_available;
   end else if(in_data_available || activation_in_progress) begin
      cycle_count = cycle_count + 1;

      for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
         if(activation_type==1'b1) begin // tanH
            slope_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= data_slope_flopped[i*8 +: 8] * inp_data_flopped[i*`DWIDTH +:`DWIDTH];
            data_intercept_flopped[i*8 +: 8] <= data_intercept[i*8 +: 8];
            data_intercept_delayed[i*8 +: 8] <= data_intercept_flopped[i*8 +: 8];
            intercept_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= slope_applied_data_internal[i*`DWIDTH +:`DWIDTH] + data_intercept_delayed[i*8 +: 8];
         end else begin // ReLU
            relu_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= inp_data[i*`DWIDTH] ? {`DWIDTH{1'b0}} : inp_data[i*`DWIDTH +:`DWIDTH];
         end
      end   

      //TANH needs 1 extra cycle
      if (activation_type==1'b1) begin
         if (cycle_count==3) begin
            out_data_available_internal <= 1;
         end
      end else begin
         if (cycle_count==2) begin
           out_data_available_internal <= 1;
         end
      end

      //TANH needs 1 extra cycle
      if (activation_type==1'b1) begin
        if(cycle_count==(`DESIGN_SIZE+2)) begin
           done_activation_internal <= 1'b1;
           activation_in_progress <= 0;
        end
        else begin
           activation_in_progress <= 1;
        end
      end else begin
        if(cycle_count==(`DESIGN_SIZE+1)) begin
           done_activation_internal <= 1'b1;
           activation_in_progress <= 0;
        end
        else begin
           activation_in_progress <= 1;
        end
      end
   end
   else begin
      slope_applied_data_internal     <= 0;
      intercept_applied_data_internal <= 0; 
      relu_applied_data_internal      <= 0; 
      data_intercept_delayed      <= 0;
      data_intercept_flopped      <= 0;
      done_activation_internal    <= 0;
      out_data_available_internal <= 0;
      cycle_count                 <= 0;
      activation_in_progress      <= 0;
   end
end

assign out_data_internal = (activation_type) ? intercept_applied_data_internal : relu_applied_data_internal;

//Our equation of tanh is Y=AX+B
//A is the slope and B is the intercept.
//We store A in one LUT and B in another.
//LUT for the slope
always @(address) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
    case (address[i*4+:4])
      4'b0000: data_slope[i*8+:8] = 8'd0;
      4'b0001: data_slope[i*8+:8] = 8'd0;
      4'b0010: data_slope[i*8+:8] = 8'd2;
      4'b0011: data_slope[i*8+:8] = 8'd3;
      4'b0100: data_slope[i*8+:8] = 8'd4;
      4'b0101: data_slope[i*8+:8] = 8'd0;
      4'b0110: data_slope[i*8+:8] = 8'd4;
      4'b0111: data_slope[i*8+:8] = 8'd3;
      4'b1000: data_slope[i*8+:8] = 8'd2;
      4'b1001: data_slope[i*8+:8] = 8'd0;
      4'b1010: data_slope[i*8+:8] = 8'd0;
      default: data_slope[i*8+:8] = 8'd0;
    endcase  
    end
end

//LUT for the intercept
always @(address) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
    case (address[i*4+:4])
      4'b0000: data_intercept[i*8+:8] = 8'd127;
      4'b0001: data_intercept[i*8+:8] = 8'd99;
      4'b0010: data_intercept[i*8+:8] = 8'd46;
      4'b0011: data_intercept[i*8+:8] = 8'd18;
      4'b0100: data_intercept[i*8+:8] = 8'd0;
      4'b0101: data_intercept[i*8+:8] = 8'd0;
      4'b0110: data_intercept[i*8+:8] = 8'd0;
      4'b0111: data_intercept[i*8+:8] = -8'd18;
      4'b1000: data_intercept[i*8+:8] = -8'd46;
      4'b1001: data_intercept[i*8+:8] = -8'd99;
      4'b1010: data_intercept[i*8+:8] = -8'd127;
      default: data_intercept[i*8+:8] = 8'd0;
    endcase  
    end
end

//Logic to find address
always @(inp_data) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
        if((inp_data[i*`DWIDTH +:`DWIDTH])>=90) begin
           address[i*4+:4] = 4'b0000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=39 && (inp_data[i*`DWIDTH +:`DWIDTH])<90) begin
           address[i*4+:4] = 4'b0001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=28 && (inp_data[i*`DWIDTH +:`DWIDTH])<39) begin
           address[i*4+:4] = 4'b0010;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=16 && (inp_data[i*`DWIDTH +:`DWIDTH])<28) begin
           address[i*4+:4] = 4'b0011;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=1 && (inp_data[i*`DWIDTH +:`DWIDTH])<16) begin
           address[i*4+:4] = 4'b0100;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])==0) begin
           address[i*4+:4] = 4'b0101;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-16 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-1) begin
           address[i*4+:4] = 4'b0110;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-28 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-16) begin
           address[i*4+:4] = 4'b0111;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-39 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-28) begin
           address[i*4+:4] = 4'b1000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-90 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-39) begin
           address[i*4+:4] = 4'b1001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])<=-90) begin
           address[i*4+:4] = 4'b1010;
        end
        else begin
           address[i*4+:4] = 4'b0101;
        end
    end
end

//Adding a dummy signal to use validity_mask input, to make ODIN happy
//TODO: Need to correctly use validity_mask
wire [`MASK_WIDTH-1:0] dummy;
assign dummy = validity_mask;

endmodule
`define DWIDTH 8
`define DESIGN_SIZE 32
`define MASK_WIDTH 2

module activation_32_8bit(
    input activation_type,
    input enable_activation,
    input in_data_available,
    input [`DESIGN_SIZE*`DWIDTH-1:0] inp_data,
    output [`DESIGN_SIZE*`DWIDTH-1:0] out_data,
    output out_data_available,
    input [`MASK_WIDTH-1:0] validity_mask,
    output done_activation,
    input clk,
    input reset
);

reg  done_activation_internal;
reg  out_data_available_internal;
wire [`DESIGN_SIZE*`DWIDTH-1:0] out_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] slope_applied_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] intercept_applied_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] relu_applied_data_internal;
reg [31:0] i;
reg [31:0] cycle_count;
reg activation_in_progress;

reg [(`DESIGN_SIZE*4)-1:0] address;
reg [(`DESIGN_SIZE*8)-1:0] data_slope;
reg [(`DESIGN_SIZE*8)-1:0] data_slope_flopped;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept_delayed;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept_flopped;

reg in_data_available_flopped;
reg [`DESIGN_SIZE*`DWIDTH-1:0] inp_data_flopped;

always @(posedge clk) begin
  if (reset) begin
    inp_data_flopped <= 0;
    data_slope_flopped <= 0;
  end else begin
    inp_data_flopped <= inp_data;
    data_slope_flopped <= data_slope;
  end
end

// If the activation block is not enabled, just forward the input data
assign out_data             = enable_activation ? out_data_internal : inp_data_flopped;
assign done_activation      = enable_activation ? done_activation_internal : 1'b1;
assign out_data_available   = enable_activation ? out_data_available_internal : in_data_available_flopped;

always @(posedge clk) begin
   if (reset || ~enable_activation) begin
      slope_applied_data_internal     <= 0;
      intercept_applied_data_internal <= 0; 
      relu_applied_data_internal      <= 0; 
      data_intercept_delayed      <= 0;
      data_intercept_flopped      <= 0;
      done_activation_internal    <= 0;
      out_data_available_internal <= 0;
      cycle_count                 <= 0;
      activation_in_progress      <= 0;
      in_data_available_flopped <= in_data_available;
   end else if(in_data_available || activation_in_progress) begin
      cycle_count = cycle_count + 1;

      for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
         if(activation_type==1'b1) begin // tanH
            slope_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= data_slope_flopped[i*8 +: 8] * inp_data_flopped[i*`DWIDTH +:`DWIDTH];
            data_intercept_flopped[i*8 +: 8] <= data_intercept[i*8 +: 8];
            data_intercept_delayed[i*8 +: 8] <= data_intercept_flopped[i*8 +: 8];
            intercept_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= slope_applied_data_internal[i*`DWIDTH +:`DWIDTH] + data_intercept_delayed[i*8 +: 8];
         end else begin // ReLU
            relu_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= inp_data[i*`DWIDTH] ? {`DWIDTH{1'b0}} : inp_data[i*`DWIDTH +:`DWIDTH];
         end
      end   

      //TANH needs 1 extra cycle
      if (activation_type==1'b1) begin
         if (cycle_count==3) begin
            out_data_available_internal <= 1;
         end
      end else begin
         if (cycle_count==2) begin
           out_data_available_internal <= 1;
         end
      end

      //TANH needs 1 extra cycle
      if (activation_type==1'b1) begin
        if(cycle_count==(`DESIGN_SIZE+2)) begin
           done_activation_internal <= 1'b1;
           activation_in_progress <= 0;
        end
        else begin
           activation_in_progress <= 1;
        end
      end else begin
        if(cycle_count==(`DESIGN_SIZE+1)) begin
           done_activation_internal <= 1'b1;
           activation_in_progress <= 0;
        end
        else begin
           activation_in_progress <= 1;
        end
      end
   end
   else begin
      slope_applied_data_internal     <= 0;
      intercept_applied_data_internal <= 0; 
      relu_applied_data_internal      <= 0; 
      data_intercept_delayed      <= 0;
      data_intercept_flopped      <= 0;
      done_activation_internal    <= 0;
      out_data_available_internal <= 0;
      cycle_count                 <= 0;
      activation_in_progress      <= 0;
   end
end

assign out_data_internal = (activation_type) ? intercept_applied_data_internal : relu_applied_data_internal;

//Our equation of tanh is Y=AX+B
//A is the slope and B is the intercept.
//We store A in one LUT and B in another.
//LUT for the slope
always @(address) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
    case (address[i*4+:4])
      4'b0000: data_slope[i*8+:8] = 8'd0;
      4'b0001: data_slope[i*8+:8] = 8'd0;
      4'b0010: data_slope[i*8+:8] = 8'd2;
      4'b0011: data_slope[i*8+:8] = 8'd3;
      4'b0100: data_slope[i*8+:8] = 8'd4;
      4'b0101: data_slope[i*8+:8] = 8'd0;
      4'b0110: data_slope[i*8+:8] = 8'd4;
      4'b0111: data_slope[i*8+:8] = 8'd3;
      4'b1000: data_slope[i*8+:8] = 8'd2;
      4'b1001: data_slope[i*8+:8] = 8'd0;
      4'b1010: data_slope[i*8+:8] = 8'd0;
      default: data_slope[i*8+:8] = 8'd0;
    endcase  
    end
end

//LUT for the intercept
always @(address) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
    case (address[i*4+:4])
      4'b0000: data_intercept[i*8+:8] = 8'd127;
      4'b0001: data_intercept[i*8+:8] = 8'd99;
      4'b0010: data_intercept[i*8+:8] = 8'd46;
      4'b0011: data_intercept[i*8+:8] = 8'd18;
      4'b0100: data_intercept[i*8+:8] = 8'd0;
      4'b0101: data_intercept[i*8+:8] = 8'd0;
      4'b0110: data_intercept[i*8+:8] = 8'd0;
      4'b0111: data_intercept[i*8+:8] = -8'd18;
      4'b1000: data_intercept[i*8+:8] = -8'd46;
      4'b1001: data_intercept[i*8+:8] = -8'd99;
      4'b1010: data_intercept[i*8+:8] = -8'd127;
      default: data_intercept[i*8+:8] = 8'd0;
    endcase  
    end
end

//Logic to find address
always @(inp_data) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
        if((inp_data[i*`DWIDTH +:`DWIDTH])>=90) begin
           address[i*4+:4] = 4'b0000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=39 && (inp_data[i*`DWIDTH +:`DWIDTH])<90) begin
           address[i*4+:4] = 4'b0001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=28 && (inp_data[i*`DWIDTH +:`DWIDTH])<39) begin
           address[i*4+:4] = 4'b0010;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=16 && (inp_data[i*`DWIDTH +:`DWIDTH])<28) begin
           address[i*4+:4] = 4'b0011;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=1 && (inp_data[i*`DWIDTH +:`DWIDTH])<16) begin
           address[i*4+:4] = 4'b0100;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])==0) begin
           address[i*4+:4] = 4'b0101;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-16 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-1) begin
           address[i*4+:4] = 4'b0110;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-28 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-16) begin
           address[i*4+:4] = 4'b0111;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-39 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-28) begin
           address[i*4+:4] = 4'b1000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-90 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-39) begin
           address[i*4+:4] = 4'b1001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])<=-90) begin
           address[i*4+:4] = 4'b1010;
        end
        else begin
           address[i*4+:4] = 4'b0101;
        end
    end
end

//Adding a dummy signal to use validity_mask input, to make ODIN happy
//TODO: Need to correctly use validity_mask
wire [`MASK_WIDTH-1:0] dummy;
assign dummy = validity_mask;

endmodule
module adder_tree_3stage_8bit (clk,reset,inp00,inp01,inp10,inp11,inp20,inp21,inp30,inp31,sum_out); 

input clk; 
input reset; 
input [7:0] inp00; 
input [7:0] inp01;
input [7:0] inp10; 
input [7:0] inp11;
input [7:0] inp20; 
input [7:0] inp21;
input [7:0] inp30; 
input [7:0] inp31;
output reg [15:0] sum_out;

reg [8:0] S_0_0; 
reg [8:0] S_0_1;
reg [8:0] S_0_2;
reg [8:0] S_0_3;

always@(posedge clk) begin 

S_0_0 <= inp00 + inp01; 
S_0_1 <= inp10 + inp11;
S_0_2 <= inp20 + inp21;
S_0_3 <= inp30 + inp31;

end 

reg [9:0] S_1_0;
reg [9:0] S_1_1;

always@(posedge clk) begin 

S_1_0 <= S_0_0 + S_0_1; 
S_1_1 <= S_0_2 + S_0_3;

end 

always@(posedge clk) begin 

if (reset == 1'b1) begin 
  sum_out <= 16'd0; 
end
else begin 
  sum_out <= S_1_0 + S_1_1; 
end

end 

endmodule 
module adder_tree_4stage_4bit(clk,reset,inp00,inp01,inp10,inp11,inp20,inp21,inp30,inp31,inp40,inp41,inp50,inp51,inp60,inp61,inp70,inp71,sum_out);

input clk;
input reset; 
input [3:0] inp00; 
input [3:0] inp01;
input [3:0] inp10; 
input [3:0] inp11;
input [3:0] inp20; 
input [3:0] inp21;
input [3:0] inp30; 
input [3:0] inp31;
input [3:0] inp40; 
input [3:0] inp41;
input [3:0] inp50; 
input [3:0] inp51;
input [3:0] inp60; 
input [3:0] inp61;
input [3:0] inp70; 
input [3:0] inp71;
output reg [7:0] sum_out;

reg [4:0] S_0_0; 
reg [4:0] S_0_1;
reg [4:0] S_0_2;
reg [4:0] S_0_3;
reg [4:0] S_0_4;
reg [4:0] S_0_5;
reg [4:0] S_0_6;
reg [4:0] S_0_7;

always@(posedge clk) begin 

S_0_0 <= inp00 + inp01; 
S_0_1 <= inp10 + inp11;
S_0_2 <= inp20 + inp21;
S_0_3 <= inp30 + inp31;
S_0_4 <= inp40 + inp41; 
S_0_5 <= inp50 + inp51;
S_0_6 <= inp60 + inp61;
S_0_7 <= inp70 + inp71;

end 

reg [5:0] S_1_0;
reg [5:0] S_1_1;
reg [5:0] S_1_2;
reg [5:0] S_1_3;

always@(posedge clk) begin 

S_1_0 <= S_0_0 + S_0_1; 
S_1_1 <= S_0_2 + S_0_3;
S_1_2 <= S_0_4 + S_0_5; 
S_1_3 <= S_0_6 + S_0_7;

end

reg [6:0] S_2_0; 
reg [6:0] S_2_1;

always@(posedge clk) begin 

S_2_0 <= S_1_0 + S_1_1; 
S_2_1 <= S_1_2 + S_1_3;

end

always@(posedge clk) begin 

if (reset == 1'b1) begin 
  sum_out <= 8'd0; 
end
else begin 
  sum_out <= S_2_0 + S_2_1; 
end

end 

endmodule 
module adder_tree_4stage_16bit(clk,reset,inp00,inp01,inp10,inp11,inp20,inp21,inp30,inp31,inp40,inp41,inp50,inp51,inp60,inp61,inp70,inp71,sum_out);

input clk;
input reset; 
input [15:0] inp00; 
input [15:0] inp01;
input [15:0] inp10; 
input [15:0] inp11;
input [15:0] inp20; 
input [15:0] inp21;
input [15:0] inp30; 
input [15:0] inp31;
input [15:0] inp40; 
input [15:0] inp41;
input [15:0] inp50; 
input [15:0] inp51;
input [15:0] inp60; 
input [15:0] inp61;
input [15:0] inp70; 
input [15:0] inp71;
output reg [31:0] sum_out;

reg [16:0] S_0_0; 
reg [16:0] S_0_1;
reg [16:0] S_0_2;
reg [16:0] S_0_3;
reg [16:0] S_0_4;
reg [16:0] S_0_5;
reg [16:0] S_0_6;
reg [16:0] S_0_7;

always@(posedge clk) begin 

S_0_0 <= inp00 + inp01; 
S_0_1 <= inp10 + inp11;
S_0_2 <= inp20 + inp21;
S_0_3 <= inp30 + inp31;
S_0_4 <= inp40 + inp41; 
S_0_5 <= inp50 + inp51;
S_0_6 <= inp60 + inp61;
S_0_7 <= inp70 + inp71;

end 

reg [17:0] S_1_0;
reg [17:0] S_1_1;
reg [17:0] S_1_2;
reg [17:0] S_1_3;

always@(posedge clk) begin 

S_1_0 <= S_0_0 + S_0_1; 
S_1_1 <= S_0_2 + S_0_3;
S_1_2 <= S_0_4 + S_0_5; 
S_1_3 <= S_0_6 + S_0_7;

end

reg [18:0] S_2_0; 
reg [18:0] S_2_1;

always@(posedge clk) begin 

S_2_0 <= S_1_0 + S_1_1; 
S_2_1 <= S_1_2 + S_1_3;

end

always@(posedge clk) begin 

if (reset == 1'b1) begin 
  sum_out <= 32'd0; 
end
else begin 
  sum_out <= S_2_0 + S_2_1; 
end

end 

endmodule 
module sigmoid(
input [15:0] x,
output [15:0] sig_out
);

reg [15:0] lut;
reg [5:0] address;

assign sig_out = lut;

always @(address)
begin

       case(address)
       6'd0: lut = 16'b0000000000101101; //sig(-4.5)
       6'd1: lut = 16'b0000000000110110; //sig(-4.3)
       6'd2: lut = 16'b0000000001000010; //sig(-4.1)
       6'd3: lut = 16'b0000000001010001; //sig(-3.9)
       6'd4:  lut = 16'b0000000001100010; //sig(-3.7)
       6'd5 :  lut = 16'b0000000001111000; //sig(-3.5)
       6'd6 :  lut= 16'b0000000010010001; //sig(-3.3)
       6'd7 :  lut= 16'b0000000010110000; //sig(-3.1)
       6'd8:  lut= 16'b0000000011010101; //sig(-2.9)
       6'd9 :  lut= 16'b0000000100000010; //sig(-2.7)
       6'd10 :  lut= 16'b0000000100110110; //sig(-2.5)
       6'd11 :  lut= 16'b0000000101110101; //sig(-2.3)
       6'd12 :  lut= 16'b0000000110111110; //sig(-2.1)
       6'd13 :  lut= 16'b0000001000010100; //sig(-1.9)
       6'd14 :  lut= 16'b0000001001111000; //sig(-1.7)
       6'd15 :  lut= 16'b0000001011101011; //sig(-1.5)
       6'd16 :  lut= 16'b0000001101101101; //sig(-1.3)
       6'd17:  lut= 16'b0000001111111110; //sig(-1.1)
       6'd18 :  lut= 16'b0000010010100000; //sig(-0.9)
       6'd19 :  lut= 16'b0000010101001111; //sig(-0.7)
       6'd20 :  lut= 16'b0000011000001010; //sig(-0.5)
       6'd21 :  lut= 16'b0000011011001111; //sig(-0.3)
       6'd22 :  lut= 16'b0000011110011001; //sig(-0.1)
       6'd23 :  lut= 16'b0000100001100110; //sig(0.1)
       6'd24 :  lut= 16'b0000100100110000; //sig(0.3)
       6'd25 :  lut= 16'b0000100111110101; //sig(0.5)
       6'd26 :  lut= 16'b0000101010110000; //sig(0.7)
       6'd27 :  lut= 16'b0000101101100000; //sig(0.9)
       6'd28 :  lut= 16'b0000110000000001; //sig(1.1)
       6'd29 :  lut= 16'b0000110010010010; //sig(1.3)
       6'd30 :  lut= 16'b0000110100010100; //sig(1.5)
       6'd31 :  lut= 16'b0000110110000111; //sig(1.7)
       6'd32 :  lut= 16'b0000110111101011; //sig(1.9)
       6'd33 :  lut= 16'b0000111001000001; //sig(2.1)
       6'd34 :  lut= 16'b0000111010001010; //sig(2.3)
       6'd35 :  lut= 16'b0000111011001001; //sig(2.5)
       6'd36 :  lut= 16'b0000111011111110; //sig(2.7)
       6'd37 :  lut= 16'b0000111100101010; //sig(2.9)
       6'd38 :  lut= 16'b0000111101001111; //sig(3.1)
       6'd39 :  lut= 16'b0000111101101110; //sig(3.3)
       6'd40 :  lut= 16'b0000111110000111; //sig(3.5)
       6'd41 :  lut= 16'b0000111110011101; //sig(3.7)
       6'd42 :  lut= 16'b0000111110101110; //sig(3.9)
       6'd43 :  lut= 16'b0000111110111101; //sig(4.1)
       6'd44 :  lut= 16'b0000111111001001; //sig(4.3)
       6'd45 :  lut= 16'b0000111111010011; //sig(4.5)
       6'd46 :  lut= 16'b0000111111011011; //sig(4.7)
       6'd47 :  lut= 16'b0000000000100100; //sig(-4.7)
       6'd48:   lut= 16'b0000000000000000; //0
       6'd49:   lut= 16'b0001000000000000; //1
       default: lut=0;
        endcase
end


always@(x)
begin

    case({x[15:12]})
        4'b1000:address = 6'd48;
        4'b1001:address = 6'd48;
        4'b1010:address = 6'd48;
        4'b1011:address = 6'd48;
        4'b1100:address = 6'd48;
        4'b1101:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // -3
                    begin
                       address = 6'd8;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address = 6'd9;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address = 6'd10;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd11;
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                        address =  6'd12;
                    end
        4'b1110:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // -2
                    begin
                        address =  6'd13;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address =  6'd14;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address = 6'd15;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd16;
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                        address =  6'd17;
                    end
        4'b1111:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333))  // -1
                    begin
                        address =  6'd18;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address =  6'd19;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address =  6'd20;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd21;                                                                                     
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                        address =  6'd22;
                    end
        4'b0000:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // 0
                    begin
                        address =  6'd23;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address =  6'd24;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address =  6'd25;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd26;
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                        address =  6'd27;
                    end
        4'b0001:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // 1
                    begin
                        address =  6'd28;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address =  6'd29;
                    end
                else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address =  6'd30;
                    end
                else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd31;
                    end
                else if(x[11:0] > 12'hccd)
                    begin
                       address =  6'd32;
                    end
        4'b0010:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333))  // 2
                    begin
                      address =  6'd33;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                      address =  6'd34;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                       address =  6'd35;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                       address =  6'd36;
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                       address =  6'd37;
                    end
        4'b0011:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // 3
                    begin
                       address =  6'd38;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                      address =  6'd39;
                    end
                else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                      address =  6'd40;
                    end
                else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                      address = 6'd41;
                    end
               else if(x[11:0] > 12'hccd)
                    begin
                       address = 6'd42;
                    end
        4'b0100:address = 6'd49;
        4'b0101:address = 6'd49;
        4'b0110:address = 6'd49;
        4'b0111:address = 6'd49;
       /* 4'b0100:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) //4
                    begin
                      address = lut[43];
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                       address = lut[44];
                    end
                else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                       address = lut[45];
                    end
                else if(x[11:0] > 12'h99a)
                    begin
                        address = lut[46];
                    end
        4'b0101: address = lut[46];
        4'b0110: address = lut[46];
        4'b0111: address = lut[46];  */
        default: address = 16'h1000;
        endcase

end

endmodule

